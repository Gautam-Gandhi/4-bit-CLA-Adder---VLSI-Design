magic
tech scmos
timestamp 1732090761
<< nwell >>
rect -26 -25 -2 14
rect 49 -16 172 23
rect 206 -1 246 24
rect 49 -36 85 -16
rect 206 -35 286 -1
rect 246 -40 286 -35
rect -19 -163 17 -124
rect 52 -163 100 -124
rect 126 -163 186 -124
rect 234 -163 306 -124
rect -19 -324 21 -299
rect -19 -358 131 -324
rect 184 -357 224 -352
rect 21 -363 131 -358
rect -153 -385 -117 -365
rect -153 -453 -30 -385
rect 144 -391 224 -357
rect 249 -380 285 -360
rect -19 -433 33 -394
rect 144 -416 184 -391
rect 203 -452 243 -447
rect -153 -473 -117 -453
rect 163 -471 243 -452
rect 249 -448 388 -380
rect 249 -468 285 -448
rect -19 -513 21 -488
rect 69 -510 117 -471
rect 123 -486 243 -471
rect 123 -510 203 -486
rect 163 -511 203 -510
rect -153 -561 -117 -541
rect -19 -547 61 -513
rect 21 -552 61 -547
rect -153 -629 -30 -561
rect -19 -622 33 -583
rect 69 -614 105 -575
rect 247 -594 283 -574
rect -153 -649 -117 -629
rect 247 -662 386 -594
rect 75 -710 135 -671
rect 185 -679 225 -674
rect 145 -715 225 -679
rect 247 -682 283 -662
rect -19 -749 21 -724
rect 145 -735 185 -715
rect -153 -798 -117 -778
rect -19 -783 61 -749
rect 145 -774 205 -735
rect 257 -765 297 -760
rect 21 -788 61 -783
rect -153 -866 -30 -798
rect -19 -858 33 -819
rect 81 -831 129 -792
rect 217 -799 297 -765
rect 217 -824 257 -799
rect -153 -886 -117 -866
rect 81 -935 117 -896
rect -153 -974 -117 -954
rect -153 -1013 -30 -974
rect 69 -1030 141 -991
rect -19 -1130 21 -1105
rect -153 -1179 -117 -1159
rect -19 -1164 61 -1130
rect 216 -1131 355 -1117
rect 21 -1169 61 -1164
rect 77 -1170 137 -1131
rect 148 -1156 355 -1131
rect 148 -1170 252 -1156
rect 216 -1176 252 -1170
rect -153 -1247 -30 -1179
rect -19 -1239 33 -1200
rect -153 -1267 -117 -1247
rect 87 -1293 135 -1253
rect 97 -1398 133 -1359
<< ntransistor >>
rect -15 -45 -13 -35
rect 96 -50 98 -30
rect 108 -50 110 -30
rect 131 -50 133 -30
rect 143 -50 145 -30
rect 159 -36 161 -26
rect 60 -64 62 -54
rect 217 -60 219 -50
rect 257 -60 259 -50
rect 273 -60 275 -50
rect -8 -200 -6 -180
rect 4 -200 6 -180
rect 63 -217 65 -187
rect 75 -217 77 -187
rect 87 -217 89 -187
rect 137 -234 139 -194
rect 149 -234 151 -194
rect 161 -234 163 -194
rect 173 -234 175 -194
rect 245 -251 247 -201
rect 257 -251 259 -201
rect 269 -251 271 -201
rect 281 -251 283 -201
rect 293 -251 295 -201
rect -142 -347 -140 -337
rect -106 -371 -104 -351
rect -94 -371 -92 -351
rect -71 -371 -69 -351
rect -59 -371 -57 -351
rect -43 -375 -41 -365
rect 155 -342 157 -332
rect 195 -342 197 -332
rect 211 -342 213 -332
rect 260 -342 262 -332
rect -8 -383 -6 -373
rect 32 -383 34 -373
rect 48 -383 50 -373
rect 71 -400 73 -380
rect 83 -400 85 -380
rect 106 -400 108 -380
rect 118 -400 120 -380
rect 296 -366 298 -346
rect 308 -366 310 -346
rect 331 -366 333 -346
rect 343 -366 345 -346
rect 359 -370 361 -360
rect 375 -370 377 -360
rect 174 -437 176 -427
rect 214 -437 216 -427
rect 230 -437 232 -427
rect -106 -487 -104 -467
rect -94 -487 -92 -467
rect -71 -487 -69 -467
rect -59 -487 -57 -467
rect -43 -473 -41 -463
rect -8 -470 -6 -450
rect 4 -470 6 -450
rect 20 -453 22 -443
rect -142 -501 -140 -491
rect -142 -523 -140 -513
rect -106 -547 -104 -527
rect -94 -547 -92 -527
rect -71 -547 -69 -527
rect -59 -547 -57 -527
rect 296 -482 298 -462
rect 308 -482 310 -462
rect 331 -482 333 -462
rect 343 -482 345 -462
rect 359 -468 361 -458
rect 375 -468 377 -458
rect 260 -496 262 -486
rect -43 -551 -41 -541
rect -8 -572 -6 -562
rect 32 -572 34 -562
rect 48 -572 50 -562
rect 80 -564 82 -534
rect 92 -564 94 -534
rect 104 -564 106 -534
rect 134 -564 136 -534
rect 146 -564 148 -534
rect 158 -564 160 -534
rect 258 -556 260 -546
rect 294 -580 296 -560
rect 306 -580 308 -560
rect 329 -580 331 -560
rect 341 -580 343 -560
rect 357 -584 359 -574
rect 373 -584 375 -574
rect -106 -663 -104 -643
rect -94 -663 -92 -643
rect -71 -663 -69 -643
rect -59 -663 -57 -643
rect -43 -649 -41 -639
rect -8 -659 -6 -639
rect 4 -659 6 -639
rect 20 -642 22 -632
rect 80 -651 82 -631
rect 92 -651 94 -631
rect 156 -664 158 -654
rect 196 -664 198 -654
rect 212 -664 214 -654
rect -142 -677 -140 -667
rect -142 -760 -140 -750
rect -106 -784 -104 -764
rect -94 -784 -92 -764
rect -71 -784 -69 -764
rect -59 -784 -57 -764
rect 294 -696 296 -676
rect 306 -696 308 -676
rect 329 -696 331 -676
rect 341 -696 343 -676
rect 357 -682 359 -672
rect 373 -682 375 -672
rect 258 -710 260 -700
rect -43 -788 -41 -778
rect 86 -781 88 -741
rect 98 -781 100 -741
rect 110 -781 112 -741
rect 122 -781 124 -741
rect 228 -750 230 -740
rect 268 -750 270 -740
rect 284 -750 286 -740
rect -8 -808 -6 -798
rect 32 -808 34 -798
rect 48 -808 50 -798
rect 156 -845 158 -805
rect 168 -845 170 -805
rect 180 -845 182 -805
rect 192 -845 194 -805
rect -106 -900 -104 -880
rect -94 -900 -92 -880
rect -71 -900 -69 -880
rect -59 -900 -57 -880
rect -43 -886 -41 -876
rect -8 -895 -6 -875
rect 4 -895 6 -875
rect 20 -878 22 -868
rect 92 -885 94 -855
rect 104 -885 106 -855
rect 116 -885 118 -855
rect -142 -914 -140 -904
rect -142 -936 -140 -926
rect -106 -960 -104 -940
rect -94 -960 -92 -940
rect -71 -960 -69 -940
rect -59 -960 -57 -940
rect -43 -964 -41 -954
rect 92 -972 94 -952
rect 104 -972 106 -952
rect 80 -1118 82 -1068
rect 92 -1118 94 -1068
rect 104 -1118 106 -1068
rect 116 -1118 118 -1068
rect 128 -1118 130 -1068
rect -142 -1141 -140 -1131
rect -106 -1165 -104 -1145
rect -94 -1165 -92 -1145
rect -71 -1165 -69 -1145
rect -59 -1165 -57 -1145
rect -43 -1169 -41 -1159
rect -8 -1189 -6 -1179
rect 32 -1189 34 -1179
rect 48 -1189 50 -1179
rect 88 -1241 90 -1201
rect 100 -1241 102 -1201
rect 112 -1241 114 -1201
rect 124 -1241 126 -1201
rect 263 -1190 265 -1170
rect 275 -1190 277 -1170
rect 298 -1190 300 -1170
rect 310 -1190 312 -1170
rect 326 -1176 328 -1166
rect 342 -1176 344 -1166
rect 227 -1204 229 -1194
rect -106 -1281 -104 -1261
rect -94 -1281 -92 -1261
rect -71 -1281 -69 -1261
rect -59 -1281 -57 -1261
rect -43 -1267 -41 -1257
rect -8 -1276 -6 -1256
rect 4 -1276 6 -1256
rect 20 -1259 22 -1249
rect 159 -1258 161 -1208
rect 171 -1258 173 -1208
rect 183 -1258 185 -1208
rect 195 -1258 197 -1208
rect 207 -1258 209 -1208
rect -142 -1295 -140 -1285
rect 98 -1347 100 -1317
rect 110 -1347 112 -1317
rect 122 -1347 124 -1317
rect 108 -1435 110 -1415
rect 120 -1435 122 -1415
<< ptransistor >>
rect -15 -19 -13 1
rect 60 -30 62 10
rect 72 -30 74 10
rect 96 -10 98 10
rect 131 -10 133 10
rect 159 -10 161 10
rect 217 -29 219 11
rect 233 -29 235 11
rect 257 -34 259 -14
rect 273 -34 275 -14
rect -8 -157 -6 -137
rect 4 -157 6 -137
rect 63 -157 65 -137
rect 75 -157 77 -137
rect 87 -157 89 -137
rect 137 -157 139 -137
rect 149 -157 151 -137
rect 161 -157 163 -137
rect 173 -157 175 -137
rect 245 -157 247 -137
rect 257 -157 259 -137
rect 269 -157 271 -137
rect 281 -157 283 -137
rect 293 -157 295 -137
rect -8 -352 -6 -312
rect 8 -352 10 -312
rect -142 -411 -140 -371
rect -130 -411 -128 -371
rect 32 -357 34 -337
rect 48 -357 50 -337
rect 71 -357 73 -337
rect 83 -357 85 -337
rect 106 -357 108 -337
rect 118 -357 120 -337
rect -106 -411 -104 -391
rect -71 -411 -69 -391
rect -43 -411 -41 -391
rect 155 -403 157 -363
rect 171 -403 173 -363
rect 195 -378 197 -358
rect 211 -378 213 -358
rect -8 -427 -6 -407
rect 4 -427 6 -407
rect 20 -427 22 -407
rect 260 -406 262 -366
rect 272 -406 274 -366
rect 296 -406 298 -386
rect 331 -406 333 -386
rect 359 -406 361 -386
rect 375 -406 377 -386
rect -142 -467 -140 -427
rect -130 -467 -128 -427
rect -106 -447 -104 -427
rect -71 -447 -69 -427
rect -43 -447 -41 -427
rect -8 -541 -6 -501
rect 8 -541 10 -501
rect 80 -504 82 -484
rect 92 -504 94 -484
rect 104 -504 106 -484
rect 134 -504 136 -484
rect 146 -504 148 -484
rect 158 -504 160 -484
rect 174 -498 176 -458
rect 190 -498 192 -458
rect 214 -473 216 -453
rect 230 -473 232 -453
rect 260 -462 262 -422
rect 272 -462 274 -422
rect 296 -442 298 -422
rect 331 -442 333 -422
rect 359 -442 361 -422
rect 375 -442 377 -422
rect -142 -587 -140 -547
rect -130 -587 -128 -547
rect 32 -546 34 -526
rect 48 -546 50 -526
rect -106 -587 -104 -567
rect -71 -587 -69 -567
rect -43 -587 -41 -567
rect -142 -643 -140 -603
rect -130 -643 -128 -603
rect -106 -623 -104 -603
rect -71 -623 -69 -603
rect -43 -623 -41 -603
rect -8 -616 -6 -596
rect 4 -616 6 -596
rect 20 -616 22 -596
rect 80 -608 82 -588
rect 92 -608 94 -588
rect 258 -620 260 -580
rect 270 -620 272 -580
rect 294 -620 296 -600
rect 329 -620 331 -600
rect 357 -620 359 -600
rect 373 -620 375 -600
rect 86 -704 88 -684
rect 98 -704 100 -684
rect 110 -704 112 -684
rect 122 -704 124 -684
rect 258 -676 260 -636
rect 270 -676 272 -636
rect 294 -656 296 -636
rect 329 -656 331 -636
rect 357 -656 359 -636
rect 373 -656 375 -636
rect -8 -777 -6 -737
rect 8 -777 10 -737
rect 156 -725 158 -685
rect 172 -725 174 -685
rect 196 -700 198 -680
rect 212 -700 214 -680
rect -142 -824 -140 -784
rect -130 -824 -128 -784
rect 32 -782 34 -762
rect 48 -782 50 -762
rect 156 -768 158 -748
rect 168 -768 170 -748
rect 180 -768 182 -748
rect 192 -768 194 -748
rect -106 -824 -104 -804
rect -71 -824 -69 -804
rect -43 -824 -41 -804
rect 92 -825 94 -805
rect 104 -825 106 -805
rect 116 -825 118 -805
rect -142 -880 -140 -840
rect -130 -880 -128 -840
rect -106 -860 -104 -840
rect -71 -860 -69 -840
rect -43 -860 -41 -840
rect -8 -852 -6 -832
rect 4 -852 6 -832
rect 20 -852 22 -832
rect 228 -811 230 -771
rect 244 -811 246 -771
rect 268 -786 270 -766
rect 284 -786 286 -766
rect 92 -929 94 -909
rect 104 -929 106 -909
rect -142 -1000 -140 -960
rect -130 -1000 -128 -960
rect -106 -1000 -104 -980
rect -71 -1000 -69 -980
rect -43 -1000 -41 -980
rect 80 -1024 82 -1004
rect 92 -1024 94 -1004
rect 104 -1024 106 -1004
rect 116 -1024 118 -1004
rect 128 -1024 130 -1004
rect -8 -1158 -6 -1118
rect 8 -1158 10 -1118
rect -142 -1205 -140 -1165
rect -130 -1205 -128 -1165
rect 32 -1163 34 -1143
rect 48 -1163 50 -1143
rect 88 -1164 90 -1144
rect 100 -1164 102 -1144
rect 112 -1164 114 -1144
rect 124 -1164 126 -1144
rect 159 -1164 161 -1144
rect 171 -1164 173 -1144
rect 183 -1164 185 -1144
rect 195 -1164 197 -1144
rect 207 -1164 209 -1144
rect -106 -1205 -104 -1185
rect -71 -1205 -69 -1185
rect -43 -1205 -41 -1185
rect -142 -1261 -140 -1221
rect -130 -1261 -128 -1221
rect -106 -1241 -104 -1221
rect -71 -1241 -69 -1221
rect -43 -1241 -41 -1221
rect -8 -1233 -6 -1213
rect 4 -1233 6 -1213
rect 20 -1233 22 -1213
rect 227 -1170 229 -1130
rect 239 -1170 241 -1130
rect 263 -1150 265 -1130
rect 298 -1150 300 -1130
rect 326 -1150 328 -1130
rect 342 -1150 344 -1130
rect 98 -1287 100 -1267
rect 110 -1287 112 -1267
rect 122 -1287 124 -1267
rect 108 -1392 110 -1372
rect 120 -1392 122 -1372
<< ndiffusion >>
rect -16 -45 -15 -35
rect -13 -45 -12 -35
rect 95 -50 96 -30
rect 98 -50 108 -30
rect 110 -50 111 -30
rect 130 -50 131 -30
rect 133 -50 143 -30
rect 145 -50 146 -30
rect 158 -36 159 -26
rect 161 -36 162 -26
rect 59 -64 60 -54
rect 62 -64 63 -54
rect 216 -60 217 -50
rect 219 -60 220 -50
rect 256 -60 257 -50
rect 259 -60 260 -50
rect 272 -60 273 -50
rect 275 -60 276 -50
rect -9 -200 -8 -180
rect -6 -200 4 -180
rect 6 -200 7 -180
rect 62 -217 63 -187
rect 65 -217 75 -187
rect 77 -217 87 -187
rect 89 -217 90 -187
rect 136 -234 137 -194
rect 139 -234 149 -194
rect 151 -234 161 -194
rect 163 -234 173 -194
rect 175 -234 176 -194
rect 244 -251 245 -201
rect 247 -251 257 -201
rect 259 -251 269 -201
rect 271 -251 281 -201
rect 283 -251 293 -201
rect 295 -251 296 -201
rect -143 -347 -142 -337
rect -140 -347 -139 -337
rect -107 -371 -106 -351
rect -104 -371 -94 -351
rect -92 -371 -91 -351
rect -72 -371 -71 -351
rect -69 -371 -59 -351
rect -57 -371 -56 -351
rect -44 -375 -43 -365
rect -41 -375 -40 -365
rect 154 -342 155 -332
rect 157 -342 158 -332
rect 194 -342 195 -332
rect 197 -342 198 -332
rect 210 -342 211 -332
rect 213 -342 214 -332
rect 259 -342 260 -332
rect 262 -342 263 -332
rect -9 -383 -8 -373
rect -6 -383 -5 -373
rect 31 -383 32 -373
rect 34 -383 35 -373
rect 47 -383 48 -373
rect 50 -383 51 -373
rect 70 -400 71 -380
rect 73 -400 83 -380
rect 85 -400 86 -380
rect 105 -400 106 -380
rect 108 -400 118 -380
rect 120 -400 121 -380
rect 295 -366 296 -346
rect 298 -366 308 -346
rect 310 -366 311 -346
rect 330 -366 331 -346
rect 333 -366 343 -346
rect 345 -366 346 -346
rect 358 -370 359 -360
rect 361 -370 362 -360
rect 374 -370 375 -360
rect 377 -370 378 -360
rect 173 -437 174 -427
rect 176 -437 177 -427
rect 213 -437 214 -427
rect 216 -437 217 -427
rect 229 -437 230 -427
rect 232 -437 233 -427
rect -107 -487 -106 -467
rect -104 -487 -94 -467
rect -92 -487 -91 -467
rect -72 -487 -71 -467
rect -69 -487 -59 -467
rect -57 -487 -56 -467
rect -44 -473 -43 -463
rect -41 -473 -40 -463
rect -9 -470 -8 -450
rect -6 -470 4 -450
rect 6 -470 7 -450
rect 19 -453 20 -443
rect 22 -453 23 -443
rect -143 -501 -142 -491
rect -140 -501 -139 -491
rect -143 -523 -142 -513
rect -140 -523 -139 -513
rect -107 -547 -106 -527
rect -104 -547 -94 -527
rect -92 -547 -91 -527
rect -72 -547 -71 -527
rect -69 -547 -59 -527
rect -57 -547 -56 -527
rect 295 -482 296 -462
rect 298 -482 308 -462
rect 310 -482 311 -462
rect 330 -482 331 -462
rect 333 -482 343 -462
rect 345 -482 346 -462
rect 358 -468 359 -458
rect 361 -468 362 -458
rect 374 -468 375 -458
rect 377 -468 378 -458
rect 259 -496 260 -486
rect 262 -496 263 -486
rect -44 -551 -43 -541
rect -41 -551 -40 -541
rect -9 -572 -8 -562
rect -6 -572 -5 -562
rect 31 -572 32 -562
rect 34 -572 35 -562
rect 47 -572 48 -562
rect 50 -572 51 -562
rect 79 -564 80 -534
rect 82 -564 92 -534
rect 94 -564 104 -534
rect 106 -564 107 -534
rect 133 -564 134 -534
rect 136 -564 146 -534
rect 148 -564 158 -534
rect 160 -564 161 -534
rect 257 -556 258 -546
rect 260 -556 261 -546
rect 293 -580 294 -560
rect 296 -580 306 -560
rect 308 -580 309 -560
rect 328 -580 329 -560
rect 331 -580 341 -560
rect 343 -580 344 -560
rect 356 -584 357 -574
rect 359 -584 360 -574
rect 372 -584 373 -574
rect 375 -584 376 -574
rect -107 -663 -106 -643
rect -104 -663 -94 -643
rect -92 -663 -91 -643
rect -72 -663 -71 -643
rect -69 -663 -59 -643
rect -57 -663 -56 -643
rect -44 -649 -43 -639
rect -41 -649 -40 -639
rect -9 -659 -8 -639
rect -6 -659 4 -639
rect 6 -659 7 -639
rect 19 -642 20 -632
rect 22 -642 23 -632
rect 79 -651 80 -631
rect 82 -651 92 -631
rect 94 -651 95 -631
rect 155 -664 156 -654
rect 158 -664 159 -654
rect 195 -664 196 -654
rect 198 -664 199 -654
rect 211 -664 212 -654
rect 214 -664 215 -654
rect -143 -677 -142 -667
rect -140 -677 -139 -667
rect -143 -760 -142 -750
rect -140 -760 -139 -750
rect -107 -784 -106 -764
rect -104 -784 -94 -764
rect -92 -784 -91 -764
rect -72 -784 -71 -764
rect -69 -784 -59 -764
rect -57 -784 -56 -764
rect 293 -696 294 -676
rect 296 -696 306 -676
rect 308 -696 309 -676
rect 328 -696 329 -676
rect 331 -696 341 -676
rect 343 -696 344 -676
rect 356 -682 357 -672
rect 359 -682 360 -672
rect 372 -682 373 -672
rect 375 -682 376 -672
rect 257 -710 258 -700
rect 260 -710 261 -700
rect -44 -788 -43 -778
rect -41 -788 -40 -778
rect 85 -781 86 -741
rect 88 -781 98 -741
rect 100 -781 110 -741
rect 112 -781 122 -741
rect 124 -781 125 -741
rect 227 -750 228 -740
rect 230 -750 231 -740
rect 267 -750 268 -740
rect 270 -750 271 -740
rect 283 -750 284 -740
rect 286 -750 287 -740
rect -9 -808 -8 -798
rect -6 -808 -5 -798
rect 31 -808 32 -798
rect 34 -808 35 -798
rect 47 -808 48 -798
rect 50 -808 51 -798
rect 155 -845 156 -805
rect 158 -845 168 -805
rect 170 -845 180 -805
rect 182 -845 192 -805
rect 194 -845 195 -805
rect -107 -900 -106 -880
rect -104 -900 -94 -880
rect -92 -900 -91 -880
rect -72 -900 -71 -880
rect -69 -900 -59 -880
rect -57 -900 -56 -880
rect -44 -886 -43 -876
rect -41 -886 -40 -876
rect -9 -895 -8 -875
rect -6 -895 4 -875
rect 6 -895 7 -875
rect 19 -878 20 -868
rect 22 -878 23 -868
rect 91 -885 92 -855
rect 94 -885 104 -855
rect 106 -885 116 -855
rect 118 -885 119 -855
rect -143 -914 -142 -904
rect -140 -914 -139 -904
rect -143 -936 -142 -926
rect -140 -936 -139 -926
rect -107 -960 -106 -940
rect -104 -960 -94 -940
rect -92 -960 -91 -940
rect -72 -960 -71 -940
rect -69 -960 -59 -940
rect -57 -960 -56 -940
rect -44 -964 -43 -954
rect -41 -964 -40 -954
rect 91 -972 92 -952
rect 94 -972 104 -952
rect 106 -972 107 -952
rect 79 -1118 80 -1068
rect 82 -1118 92 -1068
rect 94 -1118 104 -1068
rect 106 -1118 116 -1068
rect 118 -1118 128 -1068
rect 130 -1118 131 -1068
rect -143 -1141 -142 -1131
rect -140 -1141 -139 -1131
rect -107 -1165 -106 -1145
rect -104 -1165 -94 -1145
rect -92 -1165 -91 -1145
rect -72 -1165 -71 -1145
rect -69 -1165 -59 -1145
rect -57 -1165 -56 -1145
rect -44 -1169 -43 -1159
rect -41 -1169 -40 -1159
rect -9 -1189 -8 -1179
rect -6 -1189 -5 -1179
rect 31 -1189 32 -1179
rect 34 -1189 35 -1179
rect 47 -1189 48 -1179
rect 50 -1189 51 -1179
rect 87 -1241 88 -1201
rect 90 -1241 100 -1201
rect 102 -1241 112 -1201
rect 114 -1241 124 -1201
rect 126 -1241 127 -1201
rect 262 -1190 263 -1170
rect 265 -1190 275 -1170
rect 277 -1190 278 -1170
rect 297 -1190 298 -1170
rect 300 -1190 310 -1170
rect 312 -1190 313 -1170
rect 325 -1176 326 -1166
rect 328 -1176 329 -1166
rect 341 -1176 342 -1166
rect 344 -1176 345 -1166
rect 226 -1204 227 -1194
rect 229 -1204 230 -1194
rect -107 -1281 -106 -1261
rect -104 -1281 -94 -1261
rect -92 -1281 -91 -1261
rect -72 -1281 -71 -1261
rect -69 -1281 -59 -1261
rect -57 -1281 -56 -1261
rect -44 -1267 -43 -1257
rect -41 -1267 -40 -1257
rect -9 -1276 -8 -1256
rect -6 -1276 4 -1256
rect 6 -1276 7 -1256
rect 19 -1259 20 -1249
rect 22 -1259 23 -1249
rect 158 -1258 159 -1208
rect 161 -1258 171 -1208
rect 173 -1258 183 -1208
rect 185 -1258 195 -1208
rect 197 -1258 207 -1208
rect 209 -1258 210 -1208
rect -143 -1295 -142 -1285
rect -140 -1295 -139 -1285
rect 97 -1347 98 -1317
rect 100 -1347 110 -1317
rect 112 -1347 122 -1317
rect 124 -1347 125 -1317
rect 107 -1435 108 -1415
rect 110 -1435 120 -1415
rect 122 -1435 123 -1415
<< pdiffusion >>
rect -16 -19 -15 1
rect -13 -19 -12 1
rect 59 -30 60 10
rect 62 -30 72 10
rect 74 -30 75 10
rect 95 -10 96 10
rect 98 -10 99 10
rect 130 -10 131 10
rect 133 -10 134 10
rect 158 -10 159 10
rect 161 -10 162 10
rect 216 -29 217 11
rect 219 -29 220 11
rect 232 -29 233 11
rect 235 -29 236 11
rect 256 -34 257 -14
rect 259 -34 260 -14
rect 272 -34 273 -14
rect 275 -34 276 -14
rect -9 -157 -8 -137
rect -6 -157 -5 -137
rect 3 -157 4 -137
rect 6 -157 7 -137
rect 62 -157 63 -137
rect 65 -157 66 -137
rect 74 -157 75 -137
rect 77 -157 78 -137
rect 86 -157 87 -137
rect 89 -157 90 -137
rect 136 -157 137 -137
rect 139 -157 140 -137
rect 148 -157 149 -137
rect 151 -157 152 -137
rect 160 -157 161 -137
rect 163 -157 164 -137
rect 172 -157 173 -137
rect 175 -157 176 -137
rect 244 -157 245 -137
rect 247 -157 248 -137
rect 256 -157 257 -137
rect 259 -157 260 -137
rect 268 -157 269 -137
rect 271 -157 272 -137
rect 280 -157 281 -137
rect 283 -157 284 -137
rect 292 -157 293 -137
rect 295 -157 296 -137
rect -9 -352 -8 -312
rect -6 -352 -5 -312
rect 7 -352 8 -312
rect 10 -352 11 -312
rect -143 -411 -142 -371
rect -140 -411 -130 -371
rect -128 -411 -127 -371
rect 31 -357 32 -337
rect 34 -357 35 -337
rect 47 -357 48 -337
rect 50 -357 51 -337
rect 70 -357 71 -337
rect 73 -357 74 -337
rect 82 -357 83 -337
rect 85 -357 86 -337
rect 105 -357 106 -337
rect 108 -357 109 -337
rect 117 -357 118 -337
rect 120 -357 121 -337
rect -107 -411 -106 -391
rect -104 -411 -103 -391
rect -72 -411 -71 -391
rect -69 -411 -68 -391
rect -44 -411 -43 -391
rect -41 -411 -40 -391
rect 154 -403 155 -363
rect 157 -403 158 -363
rect 170 -403 171 -363
rect 173 -403 174 -363
rect 194 -378 195 -358
rect 197 -378 198 -358
rect 210 -378 211 -358
rect 213 -378 214 -358
rect -9 -427 -8 -407
rect -6 -427 -5 -407
rect 3 -427 4 -407
rect 6 -427 7 -407
rect 19 -427 20 -407
rect 22 -427 23 -407
rect 259 -406 260 -366
rect 262 -406 272 -366
rect 274 -406 275 -366
rect 295 -406 296 -386
rect 298 -406 299 -386
rect 330 -406 331 -386
rect 333 -406 334 -386
rect 358 -406 359 -386
rect 361 -406 362 -386
rect 374 -406 375 -386
rect 377 -406 378 -386
rect -143 -467 -142 -427
rect -140 -467 -130 -427
rect -128 -467 -127 -427
rect -107 -447 -106 -427
rect -104 -447 -103 -427
rect -72 -447 -71 -427
rect -69 -447 -68 -427
rect -44 -447 -43 -427
rect -41 -447 -40 -427
rect -9 -541 -8 -501
rect -6 -541 -5 -501
rect 7 -541 8 -501
rect 10 -541 11 -501
rect 79 -504 80 -484
rect 82 -504 83 -484
rect 91 -504 92 -484
rect 94 -504 95 -484
rect 103 -504 104 -484
rect 106 -504 107 -484
rect 133 -504 134 -484
rect 136 -504 137 -484
rect 145 -504 146 -484
rect 148 -504 149 -484
rect 157 -504 158 -484
rect 160 -504 161 -484
rect 173 -498 174 -458
rect 176 -498 177 -458
rect 189 -498 190 -458
rect 192 -498 193 -458
rect 213 -473 214 -453
rect 216 -473 217 -453
rect 229 -473 230 -453
rect 232 -473 233 -453
rect 259 -462 260 -422
rect 262 -462 272 -422
rect 274 -462 275 -422
rect 295 -442 296 -422
rect 298 -442 299 -422
rect 330 -442 331 -422
rect 333 -442 334 -422
rect 358 -442 359 -422
rect 361 -442 362 -422
rect 374 -442 375 -422
rect 377 -442 378 -422
rect -143 -587 -142 -547
rect -140 -587 -130 -547
rect -128 -587 -127 -547
rect 31 -546 32 -526
rect 34 -546 35 -526
rect 47 -546 48 -526
rect 50 -546 51 -526
rect -107 -587 -106 -567
rect -104 -587 -103 -567
rect -72 -587 -71 -567
rect -69 -587 -68 -567
rect -44 -587 -43 -567
rect -41 -587 -40 -567
rect -143 -643 -142 -603
rect -140 -643 -130 -603
rect -128 -643 -127 -603
rect -107 -623 -106 -603
rect -104 -623 -103 -603
rect -72 -623 -71 -603
rect -69 -623 -68 -603
rect -44 -623 -43 -603
rect -41 -623 -40 -603
rect -9 -616 -8 -596
rect -6 -616 -5 -596
rect 3 -616 4 -596
rect 6 -616 7 -596
rect 19 -616 20 -596
rect 22 -616 23 -596
rect 79 -608 80 -588
rect 82 -608 83 -588
rect 91 -608 92 -588
rect 94 -608 95 -588
rect 257 -620 258 -580
rect 260 -620 270 -580
rect 272 -620 273 -580
rect 293 -620 294 -600
rect 296 -620 297 -600
rect 328 -620 329 -600
rect 331 -620 332 -600
rect 356 -620 357 -600
rect 359 -620 360 -600
rect 372 -620 373 -600
rect 375 -620 376 -600
rect 85 -704 86 -684
rect 88 -704 89 -684
rect 97 -704 98 -684
rect 100 -704 101 -684
rect 109 -704 110 -684
rect 112 -704 113 -684
rect 121 -704 122 -684
rect 124 -704 125 -684
rect 257 -676 258 -636
rect 260 -676 270 -636
rect 272 -676 273 -636
rect 293 -656 294 -636
rect 296 -656 297 -636
rect 328 -656 329 -636
rect 331 -656 332 -636
rect 356 -656 357 -636
rect 359 -656 360 -636
rect 372 -656 373 -636
rect 375 -656 376 -636
rect -9 -777 -8 -737
rect -6 -777 -5 -737
rect 7 -777 8 -737
rect 10 -777 11 -737
rect 155 -725 156 -685
rect 158 -725 159 -685
rect 171 -725 172 -685
rect 174 -725 175 -685
rect 195 -700 196 -680
rect 198 -700 199 -680
rect 211 -700 212 -680
rect 214 -700 215 -680
rect -143 -824 -142 -784
rect -140 -824 -130 -784
rect -128 -824 -127 -784
rect 31 -782 32 -762
rect 34 -782 35 -762
rect 47 -782 48 -762
rect 50 -782 51 -762
rect 155 -768 156 -748
rect 158 -768 159 -748
rect 167 -768 168 -748
rect 170 -768 171 -748
rect 179 -768 180 -748
rect 182 -768 183 -748
rect 191 -768 192 -748
rect 194 -768 195 -748
rect -107 -824 -106 -804
rect -104 -824 -103 -804
rect -72 -824 -71 -804
rect -69 -824 -68 -804
rect -44 -824 -43 -804
rect -41 -824 -40 -804
rect 91 -825 92 -805
rect 94 -825 95 -805
rect 103 -825 104 -805
rect 106 -825 107 -805
rect 115 -825 116 -805
rect 118 -825 119 -805
rect -143 -880 -142 -840
rect -140 -880 -130 -840
rect -128 -880 -127 -840
rect -107 -860 -106 -840
rect -104 -860 -103 -840
rect -72 -860 -71 -840
rect -69 -860 -68 -840
rect -44 -860 -43 -840
rect -41 -860 -40 -840
rect -9 -852 -8 -832
rect -6 -852 -5 -832
rect 3 -852 4 -832
rect 6 -852 7 -832
rect 19 -852 20 -832
rect 22 -852 23 -832
rect 227 -811 228 -771
rect 230 -811 231 -771
rect 243 -811 244 -771
rect 246 -811 247 -771
rect 267 -786 268 -766
rect 270 -786 271 -766
rect 283 -786 284 -766
rect 286 -786 287 -766
rect 91 -929 92 -909
rect 94 -929 95 -909
rect 103 -929 104 -909
rect 106 -929 107 -909
rect -143 -1000 -142 -960
rect -140 -1000 -130 -960
rect -128 -1000 -127 -960
rect -107 -1000 -106 -980
rect -104 -1000 -103 -980
rect -72 -1000 -71 -980
rect -69 -1000 -68 -980
rect -44 -1000 -43 -980
rect -41 -1000 -40 -980
rect 79 -1024 80 -1004
rect 82 -1024 83 -1004
rect 91 -1024 92 -1004
rect 94 -1024 95 -1004
rect 103 -1024 104 -1004
rect 106 -1024 107 -1004
rect 115 -1024 116 -1004
rect 118 -1024 119 -1004
rect 127 -1024 128 -1004
rect 130 -1024 131 -1004
rect -9 -1158 -8 -1118
rect -6 -1158 -5 -1118
rect 7 -1158 8 -1118
rect 10 -1158 11 -1118
rect -143 -1205 -142 -1165
rect -140 -1205 -130 -1165
rect -128 -1205 -127 -1165
rect 31 -1163 32 -1143
rect 34 -1163 35 -1143
rect 47 -1163 48 -1143
rect 50 -1163 51 -1143
rect 87 -1164 88 -1144
rect 90 -1164 91 -1144
rect 99 -1164 100 -1144
rect 102 -1164 103 -1144
rect 111 -1164 112 -1144
rect 114 -1164 115 -1144
rect 123 -1164 124 -1144
rect 126 -1164 127 -1144
rect 158 -1164 159 -1144
rect 161 -1164 162 -1144
rect 170 -1164 171 -1144
rect 173 -1164 174 -1144
rect 182 -1164 183 -1144
rect 185 -1164 186 -1144
rect 194 -1164 195 -1144
rect 197 -1164 198 -1144
rect 206 -1164 207 -1144
rect 209 -1164 210 -1144
rect -107 -1205 -106 -1185
rect -104 -1205 -103 -1185
rect -72 -1205 -71 -1185
rect -69 -1205 -68 -1185
rect -44 -1205 -43 -1185
rect -41 -1205 -40 -1185
rect -143 -1261 -142 -1221
rect -140 -1261 -130 -1221
rect -128 -1261 -127 -1221
rect -107 -1241 -106 -1221
rect -104 -1241 -103 -1221
rect -72 -1241 -71 -1221
rect -69 -1241 -68 -1221
rect -44 -1241 -43 -1221
rect -41 -1241 -40 -1221
rect -9 -1233 -8 -1213
rect -6 -1233 -5 -1213
rect 3 -1233 4 -1213
rect 6 -1233 7 -1213
rect 19 -1233 20 -1213
rect 22 -1233 23 -1213
rect 226 -1170 227 -1130
rect 229 -1170 239 -1130
rect 241 -1170 242 -1130
rect 262 -1150 263 -1130
rect 265 -1150 266 -1130
rect 297 -1150 298 -1130
rect 300 -1150 301 -1130
rect 325 -1150 326 -1130
rect 328 -1150 329 -1130
rect 341 -1150 342 -1130
rect 344 -1150 345 -1130
rect 97 -1287 98 -1267
rect 100 -1287 101 -1267
rect 109 -1287 110 -1267
rect 112 -1287 113 -1267
rect 121 -1287 122 -1267
rect 124 -1287 125 -1267
rect 107 -1392 108 -1372
rect 110 -1392 111 -1372
rect 119 -1392 120 -1372
rect 122 -1392 123 -1372
<< ndcontact >>
rect -20 -45 -16 -35
rect -12 -45 -8 -35
rect 91 -50 95 -30
rect 111 -50 115 -30
rect 126 -50 130 -30
rect 146 -50 150 -30
rect 154 -36 158 -26
rect 162 -36 166 -26
rect 55 -64 59 -54
rect 63 -64 67 -54
rect 212 -60 216 -50
rect 220 -60 224 -50
rect 252 -60 256 -50
rect 260 -60 264 -50
rect 268 -60 272 -50
rect 276 -60 280 -50
rect -13 -200 -9 -180
rect 7 -200 11 -180
rect 58 -217 62 -187
rect 90 -217 94 -187
rect 132 -234 136 -194
rect 176 -234 180 -194
rect 240 -251 244 -201
rect 296 -251 300 -201
rect -147 -347 -143 -337
rect -139 -347 -135 -337
rect -111 -371 -107 -351
rect -91 -371 -87 -351
rect -76 -371 -72 -351
rect -56 -371 -52 -351
rect -48 -375 -44 -365
rect -40 -375 -36 -365
rect 150 -342 154 -332
rect 158 -342 162 -332
rect 190 -342 194 -332
rect 198 -342 202 -332
rect 206 -342 210 -332
rect 214 -342 218 -332
rect 255 -342 259 -332
rect 263 -342 267 -332
rect -13 -383 -9 -373
rect -5 -383 -1 -373
rect 27 -383 31 -373
rect 35 -383 39 -373
rect 43 -383 47 -373
rect 51 -383 55 -373
rect 66 -400 70 -380
rect 86 -400 90 -380
rect 101 -400 105 -380
rect 121 -400 125 -380
rect 291 -366 295 -346
rect 311 -366 315 -346
rect 326 -366 330 -346
rect 346 -366 350 -346
rect 354 -370 358 -360
rect 362 -370 366 -360
rect 370 -370 374 -360
rect 378 -370 382 -360
rect 169 -437 173 -427
rect 177 -437 181 -427
rect 209 -437 213 -427
rect 217 -437 221 -427
rect 225 -437 229 -427
rect 233 -437 237 -427
rect -111 -487 -107 -467
rect -91 -487 -87 -467
rect -76 -487 -72 -467
rect -56 -487 -52 -467
rect -48 -473 -44 -463
rect -40 -473 -36 -463
rect -13 -470 -9 -450
rect 7 -470 11 -450
rect 15 -453 19 -443
rect 23 -453 27 -443
rect -147 -501 -143 -491
rect -139 -501 -135 -491
rect -147 -523 -143 -513
rect -139 -523 -135 -513
rect -111 -547 -107 -527
rect -91 -547 -87 -527
rect -76 -547 -72 -527
rect -56 -547 -52 -527
rect 291 -482 295 -462
rect 311 -482 315 -462
rect 326 -482 330 -462
rect 346 -482 350 -462
rect 354 -468 358 -458
rect 362 -468 366 -458
rect 370 -468 374 -458
rect 378 -468 382 -458
rect 255 -496 259 -486
rect 263 -496 267 -486
rect -48 -551 -44 -541
rect -40 -551 -36 -541
rect -13 -572 -9 -562
rect -5 -572 -1 -562
rect 27 -572 31 -562
rect 35 -572 39 -562
rect 43 -572 47 -562
rect 51 -572 55 -562
rect 75 -564 79 -534
rect 107 -564 111 -534
rect 129 -564 133 -534
rect 161 -564 165 -534
rect 253 -556 257 -546
rect 261 -556 265 -546
rect 289 -580 293 -560
rect 309 -580 313 -560
rect 324 -580 328 -560
rect 344 -580 348 -560
rect 352 -584 356 -574
rect 360 -584 364 -574
rect 368 -584 372 -574
rect 376 -584 380 -574
rect -111 -663 -107 -643
rect -91 -663 -87 -643
rect -76 -663 -72 -643
rect -56 -663 -52 -643
rect -48 -649 -44 -639
rect -40 -649 -36 -639
rect -13 -659 -9 -639
rect 7 -659 11 -639
rect 15 -642 19 -632
rect 23 -642 27 -632
rect 75 -651 79 -631
rect 95 -651 99 -631
rect 151 -664 155 -654
rect 159 -664 163 -654
rect 191 -664 195 -654
rect 199 -664 203 -654
rect 207 -664 211 -654
rect 215 -664 219 -654
rect -147 -677 -143 -667
rect -139 -677 -135 -667
rect -147 -760 -143 -750
rect -139 -760 -135 -750
rect -111 -784 -107 -764
rect -91 -784 -87 -764
rect -76 -784 -72 -764
rect -56 -784 -52 -764
rect 289 -696 293 -676
rect 309 -696 313 -676
rect 324 -696 328 -676
rect 344 -696 348 -676
rect 352 -682 356 -672
rect 360 -682 364 -672
rect 368 -682 372 -672
rect 376 -682 380 -672
rect 253 -710 257 -700
rect 261 -710 265 -700
rect -48 -788 -44 -778
rect -40 -788 -36 -778
rect 81 -781 85 -741
rect 125 -781 129 -741
rect 223 -750 227 -740
rect 231 -750 235 -740
rect 263 -750 267 -740
rect 271 -750 275 -740
rect 279 -750 283 -740
rect 287 -750 291 -740
rect -13 -808 -9 -798
rect -5 -808 -1 -798
rect 27 -808 31 -798
rect 35 -808 39 -798
rect 43 -808 47 -798
rect 51 -808 55 -798
rect 151 -845 155 -805
rect 195 -845 199 -805
rect -111 -900 -107 -880
rect -91 -900 -87 -880
rect -76 -900 -72 -880
rect -56 -900 -52 -880
rect -48 -886 -44 -876
rect -40 -886 -36 -876
rect -13 -895 -9 -875
rect 7 -895 11 -875
rect 15 -878 19 -868
rect 23 -878 27 -868
rect 87 -885 91 -855
rect 119 -885 123 -855
rect -147 -914 -143 -904
rect -139 -914 -135 -904
rect -147 -936 -143 -926
rect -139 -936 -135 -926
rect -111 -960 -107 -940
rect -91 -960 -87 -940
rect -76 -960 -72 -940
rect -56 -960 -52 -940
rect -48 -964 -44 -954
rect -40 -964 -36 -954
rect 87 -972 91 -952
rect 107 -972 111 -952
rect 75 -1118 79 -1068
rect 131 -1118 135 -1068
rect -147 -1141 -143 -1131
rect -139 -1141 -135 -1131
rect -111 -1165 -107 -1145
rect -91 -1165 -87 -1145
rect -76 -1165 -72 -1145
rect -56 -1165 -52 -1145
rect -48 -1169 -44 -1159
rect -40 -1169 -36 -1159
rect -13 -1189 -9 -1179
rect -5 -1189 -1 -1179
rect 27 -1189 31 -1179
rect 35 -1189 39 -1179
rect 43 -1189 47 -1179
rect 51 -1189 55 -1179
rect 83 -1241 87 -1201
rect 127 -1241 131 -1201
rect 258 -1190 262 -1170
rect 278 -1190 282 -1170
rect 293 -1190 297 -1170
rect 313 -1190 317 -1170
rect 321 -1176 325 -1166
rect 329 -1176 333 -1166
rect 337 -1176 341 -1166
rect 345 -1176 349 -1166
rect 222 -1204 226 -1194
rect 230 -1204 234 -1194
rect -111 -1281 -107 -1261
rect -91 -1281 -87 -1261
rect -76 -1281 -72 -1261
rect -56 -1281 -52 -1261
rect -48 -1267 -44 -1257
rect -40 -1267 -36 -1257
rect -13 -1276 -9 -1256
rect 7 -1276 11 -1256
rect 15 -1259 19 -1249
rect 23 -1259 27 -1249
rect 154 -1258 158 -1208
rect 210 -1258 214 -1208
rect -147 -1295 -143 -1285
rect -139 -1295 -135 -1285
rect 93 -1347 97 -1317
rect 125 -1347 129 -1317
rect 103 -1435 107 -1415
rect 123 -1435 127 -1415
<< pdcontact >>
rect -20 -19 -16 1
rect -12 -19 -8 1
rect 55 -30 59 10
rect 75 -30 79 10
rect 91 -10 95 10
rect 99 -10 103 10
rect 126 -10 130 10
rect 134 -10 138 10
rect 154 -10 158 10
rect 162 -10 166 10
rect 212 -29 216 11
rect 220 -29 224 11
rect 228 -29 232 11
rect 236 -29 240 11
rect 252 -34 256 -14
rect 260 -34 264 -14
rect 268 -34 272 -14
rect 276 -34 280 -14
rect -13 -157 -9 -137
rect -5 -157 3 -137
rect 7 -157 11 -137
rect 58 -157 62 -137
rect 66 -157 74 -137
rect 78 -157 86 -137
rect 90 -157 94 -137
rect 132 -157 136 -137
rect 140 -157 148 -137
rect 152 -157 160 -137
rect 164 -157 172 -137
rect 176 -157 180 -137
rect 240 -157 244 -137
rect 248 -157 256 -137
rect 260 -157 268 -137
rect 272 -157 280 -137
rect 284 -157 292 -137
rect 296 -157 300 -137
rect -13 -352 -9 -312
rect -5 -352 -1 -312
rect 3 -352 7 -312
rect 11 -352 15 -312
rect -147 -411 -143 -371
rect -127 -411 -123 -371
rect 27 -357 31 -337
rect 35 -357 39 -337
rect 43 -357 47 -337
rect 51 -357 55 -337
rect 66 -357 70 -337
rect 74 -357 82 -337
rect 86 -357 90 -337
rect 101 -357 105 -337
rect 109 -357 117 -337
rect 121 -357 125 -337
rect -111 -411 -107 -391
rect -103 -411 -99 -391
rect -76 -411 -72 -391
rect -68 -411 -64 -391
rect -48 -411 -44 -391
rect -40 -411 -36 -391
rect 150 -403 154 -363
rect 158 -403 162 -363
rect 166 -403 170 -363
rect 174 -403 178 -363
rect 190 -378 194 -358
rect 198 -378 202 -358
rect 206 -378 210 -358
rect 214 -378 218 -358
rect -13 -427 -9 -407
rect -5 -427 3 -407
rect 7 -427 11 -407
rect 15 -427 19 -407
rect 23 -427 27 -407
rect 255 -406 259 -366
rect 275 -406 279 -366
rect 291 -406 295 -386
rect 299 -406 303 -386
rect 326 -406 330 -386
rect 334 -406 338 -386
rect 354 -406 358 -386
rect 362 -406 366 -386
rect 370 -406 374 -386
rect 378 -406 382 -386
rect -147 -467 -143 -427
rect -127 -467 -123 -427
rect -111 -447 -107 -427
rect -103 -447 -99 -427
rect -76 -447 -72 -427
rect -68 -447 -64 -427
rect -48 -447 -44 -427
rect -40 -447 -36 -427
rect -13 -541 -9 -501
rect -5 -541 -1 -501
rect 3 -541 7 -501
rect 11 -541 15 -501
rect 75 -504 79 -484
rect 83 -504 91 -484
rect 95 -504 103 -484
rect 107 -504 111 -484
rect 129 -504 133 -484
rect 137 -504 145 -484
rect 149 -504 157 -484
rect 161 -504 165 -484
rect 169 -498 173 -458
rect 177 -498 181 -458
rect 185 -498 189 -458
rect 193 -498 197 -458
rect 209 -473 213 -453
rect 217 -473 221 -453
rect 225 -473 229 -453
rect 233 -473 237 -453
rect 255 -462 259 -422
rect 275 -462 279 -422
rect 291 -442 295 -422
rect 299 -442 303 -422
rect 326 -442 330 -422
rect 334 -442 338 -422
rect 354 -442 358 -422
rect 362 -442 366 -422
rect 370 -442 374 -422
rect 378 -442 382 -422
rect -147 -587 -143 -547
rect -127 -587 -123 -547
rect 27 -546 31 -526
rect 35 -546 39 -526
rect 43 -546 47 -526
rect 51 -546 55 -526
rect -111 -587 -107 -567
rect -103 -587 -99 -567
rect -76 -587 -72 -567
rect -68 -587 -64 -567
rect -48 -587 -44 -567
rect -40 -587 -36 -567
rect -147 -643 -143 -603
rect -127 -643 -123 -603
rect -111 -623 -107 -603
rect -103 -623 -99 -603
rect -76 -623 -72 -603
rect -68 -623 -64 -603
rect -48 -623 -44 -603
rect -40 -623 -36 -603
rect -13 -616 -9 -596
rect -5 -616 3 -596
rect 7 -616 11 -596
rect 15 -616 19 -596
rect 23 -616 27 -596
rect 75 -608 79 -588
rect 83 -608 91 -588
rect 95 -608 99 -588
rect 253 -620 257 -580
rect 273 -620 277 -580
rect 289 -620 293 -600
rect 297 -620 301 -600
rect 324 -620 328 -600
rect 332 -620 336 -600
rect 352 -620 356 -600
rect 360 -620 364 -600
rect 368 -620 372 -600
rect 376 -620 380 -600
rect 81 -704 85 -684
rect 89 -704 97 -684
rect 101 -704 109 -684
rect 113 -704 121 -684
rect 125 -704 129 -684
rect 253 -676 257 -636
rect 273 -676 277 -636
rect 289 -656 293 -636
rect 297 -656 301 -636
rect 324 -656 328 -636
rect 332 -656 336 -636
rect 352 -656 356 -636
rect 360 -656 364 -636
rect 368 -656 372 -636
rect 376 -656 380 -636
rect -13 -777 -9 -737
rect -5 -777 -1 -737
rect 3 -777 7 -737
rect 11 -777 15 -737
rect 151 -725 155 -685
rect 159 -725 163 -685
rect 167 -725 171 -685
rect 175 -725 179 -685
rect 191 -700 195 -680
rect 199 -700 203 -680
rect 207 -700 211 -680
rect 215 -700 219 -680
rect -147 -824 -143 -784
rect -127 -824 -123 -784
rect 27 -782 31 -762
rect 35 -782 39 -762
rect 43 -782 47 -762
rect 51 -782 55 -762
rect 151 -768 155 -748
rect 159 -768 167 -748
rect 171 -768 179 -748
rect 183 -768 191 -748
rect 195 -768 199 -748
rect -111 -824 -107 -804
rect -103 -824 -99 -804
rect -76 -824 -72 -804
rect -68 -824 -64 -804
rect -48 -824 -44 -804
rect -40 -824 -36 -804
rect 87 -825 91 -805
rect 95 -825 103 -805
rect 107 -825 115 -805
rect 119 -825 123 -805
rect -147 -880 -143 -840
rect -127 -880 -123 -840
rect -111 -860 -107 -840
rect -103 -860 -99 -840
rect -76 -860 -72 -840
rect -68 -860 -64 -840
rect -48 -860 -44 -840
rect -40 -860 -36 -840
rect -13 -852 -9 -832
rect -5 -852 3 -832
rect 7 -852 11 -832
rect 15 -852 19 -832
rect 23 -852 27 -832
rect 223 -811 227 -771
rect 231 -811 235 -771
rect 239 -811 243 -771
rect 247 -811 251 -771
rect 263 -786 267 -766
rect 271 -786 275 -766
rect 279 -786 283 -766
rect 287 -786 291 -766
rect 87 -929 91 -909
rect 95 -929 103 -909
rect 107 -929 111 -909
rect -147 -1000 -143 -960
rect -127 -1000 -123 -960
rect -111 -1000 -107 -980
rect -103 -1000 -99 -980
rect -76 -1000 -72 -980
rect -68 -1000 -64 -980
rect -48 -1000 -44 -980
rect -40 -1000 -36 -980
rect 75 -1024 79 -1004
rect 83 -1024 91 -1004
rect 95 -1024 103 -1004
rect 107 -1024 115 -1004
rect 119 -1024 127 -1004
rect 131 -1024 135 -1004
rect -13 -1158 -9 -1118
rect -5 -1158 -1 -1118
rect 3 -1158 7 -1118
rect 11 -1158 15 -1118
rect -147 -1205 -143 -1165
rect -127 -1205 -123 -1165
rect 27 -1163 31 -1143
rect 35 -1163 39 -1143
rect 43 -1163 47 -1143
rect 51 -1163 55 -1143
rect 83 -1164 87 -1144
rect 91 -1164 99 -1144
rect 103 -1164 111 -1144
rect 115 -1164 123 -1144
rect 127 -1164 131 -1144
rect 154 -1164 158 -1144
rect 162 -1164 170 -1144
rect 174 -1164 182 -1144
rect 186 -1164 194 -1144
rect 198 -1164 206 -1144
rect 210 -1164 214 -1144
rect -111 -1205 -107 -1185
rect -103 -1205 -99 -1185
rect -76 -1205 -72 -1185
rect -68 -1205 -64 -1185
rect -48 -1205 -44 -1185
rect -40 -1205 -36 -1185
rect -147 -1261 -143 -1221
rect -127 -1261 -123 -1221
rect -111 -1241 -107 -1221
rect -103 -1241 -99 -1221
rect -76 -1241 -72 -1221
rect -68 -1241 -64 -1221
rect -48 -1241 -44 -1221
rect -40 -1241 -36 -1221
rect -13 -1233 -9 -1213
rect -5 -1233 3 -1213
rect 7 -1233 11 -1213
rect 15 -1233 19 -1213
rect 23 -1233 27 -1213
rect 222 -1170 226 -1130
rect 242 -1170 246 -1130
rect 258 -1150 262 -1130
rect 266 -1150 270 -1130
rect 293 -1150 297 -1130
rect 301 -1150 305 -1130
rect 321 -1150 325 -1130
rect 329 -1150 333 -1130
rect 337 -1150 341 -1130
rect 345 -1150 349 -1130
rect 93 -1287 97 -1267
rect 101 -1287 109 -1267
rect 113 -1287 121 -1267
rect 125 -1287 129 -1267
rect 103 -1392 107 -1372
rect 111 -1392 119 -1372
rect 123 -1392 127 -1372
<< psubstratepcontact >>
rect -20 -53 -16 -49
rect -12 -53 -8 -49
rect 154 -44 158 -40
rect 162 -44 166 -40
rect 91 -58 95 -54
rect 101 -58 105 -54
rect 126 -58 130 -54
rect 136 -58 140 -54
rect 146 -58 150 -54
rect 212 -68 216 -64
rect 220 -68 224 -64
rect 252 -68 256 -64
rect 260 -68 264 -64
rect 268 -68 272 -64
rect 276 -68 280 -64
rect 55 -72 59 -68
rect 63 -72 67 -68
rect -13 -208 -9 -204
rect -3 -208 1 -204
rect 7 -208 11 -204
rect 58 -225 62 -221
rect 69 -225 73 -221
rect 79 -225 83 -221
rect 90 -225 94 -221
rect 132 -242 136 -238
rect 142 -242 146 -238
rect 154 -242 158 -238
rect 166 -242 170 -238
rect 176 -242 180 -238
rect 240 -259 244 -255
rect 250 -259 254 -255
rect 262 -259 266 -255
rect 274 -259 278 -255
rect 286 -259 290 -255
rect 296 -259 300 -255
rect -147 -333 -143 -329
rect -139 -333 -135 -329
rect -111 -347 -107 -343
rect -101 -347 -97 -343
rect -91 -347 -87 -343
rect -76 -347 -72 -343
rect -66 -347 -62 -343
rect -56 -347 -52 -343
rect 150 -328 154 -324
rect 158 -328 162 -324
rect 190 -328 194 -324
rect 198 -328 202 -324
rect 206 -328 210 -324
rect 214 -328 218 -324
rect 255 -328 259 -324
rect 263 -328 267 -324
rect -48 -361 -44 -357
rect -40 -361 -36 -357
rect 291 -342 295 -338
rect 301 -342 305 -338
rect 311 -342 315 -338
rect 326 -342 330 -338
rect 336 -342 340 -338
rect 346 -342 350 -338
rect -13 -391 -9 -387
rect -5 -391 -1 -387
rect 27 -391 31 -387
rect 35 -391 39 -387
rect 43 -391 47 -387
rect 51 -391 55 -387
rect 354 -356 358 -352
rect 362 -356 366 -352
rect 370 -356 374 -352
rect 378 -356 382 -352
rect 66 -408 70 -404
rect 76 -408 80 -404
rect 86 -408 90 -404
rect 101 -408 105 -404
rect 111 -408 115 -404
rect 121 -408 125 -404
rect 169 -423 173 -419
rect 177 -423 181 -419
rect 209 -423 213 -419
rect 217 -423 221 -419
rect 225 -423 229 -419
rect 233 -423 237 -419
rect 15 -461 19 -457
rect 25 -461 29 -457
rect -48 -481 -44 -477
rect -40 -481 -36 -477
rect -13 -478 -9 -474
rect -3 -478 1 -474
rect 7 -478 11 -474
rect -111 -495 -107 -491
rect -101 -495 -97 -491
rect -91 -495 -87 -491
rect -76 -495 -72 -491
rect -66 -495 -62 -491
rect -56 -495 -52 -491
rect -147 -509 -143 -505
rect -139 -509 -135 -505
rect -111 -523 -107 -519
rect -101 -523 -97 -519
rect -91 -523 -87 -519
rect -76 -523 -72 -519
rect -66 -523 -62 -519
rect -56 -523 -52 -519
rect -48 -537 -44 -533
rect -40 -537 -36 -533
rect 354 -476 358 -472
rect 362 -476 366 -472
rect 370 -476 374 -472
rect 378 -476 382 -472
rect 291 -490 295 -486
rect 301 -490 305 -486
rect 311 -490 315 -486
rect 326 -490 330 -486
rect 336 -490 340 -486
rect 346 -490 350 -486
rect 255 -504 259 -500
rect 263 -504 267 -500
rect 253 -542 257 -538
rect 261 -542 265 -538
rect 289 -556 293 -552
rect 299 -556 303 -552
rect 309 -556 313 -552
rect 324 -556 328 -552
rect 334 -556 338 -552
rect 344 -556 348 -552
rect 75 -572 79 -568
rect 85 -572 89 -568
rect 97 -572 101 -568
rect 107 -572 111 -568
rect 129 -572 133 -568
rect 139 -572 143 -568
rect 151 -572 155 -568
rect 161 -572 165 -568
rect -13 -580 -9 -576
rect -5 -580 -1 -576
rect 27 -580 31 -576
rect 35 -580 39 -576
rect 43 -580 47 -576
rect 352 -570 356 -566
rect 360 -570 364 -566
rect 368 -570 372 -566
rect 376 -570 380 -566
rect -48 -657 -44 -653
rect -40 -657 -36 -653
rect 15 -650 19 -646
rect 25 -650 29 -646
rect 151 -650 155 -646
rect 159 -650 163 -646
rect 191 -650 195 -646
rect 199 -650 203 -646
rect 207 -650 211 -646
rect 215 -650 219 -646
rect 75 -659 79 -655
rect 85 -659 89 -655
rect 95 -659 99 -655
rect -13 -667 -9 -663
rect -3 -667 1 -663
rect 7 -667 11 -663
rect -111 -671 -107 -667
rect -101 -671 -97 -667
rect -91 -671 -87 -667
rect -76 -671 -72 -667
rect -66 -671 -62 -667
rect -56 -671 -52 -667
rect -147 -685 -143 -681
rect -139 -685 -135 -681
rect -147 -746 -143 -742
rect -139 -746 -135 -742
rect -111 -760 -107 -756
rect -101 -760 -97 -756
rect -91 -760 -87 -756
rect -76 -760 -72 -756
rect -66 -760 -62 -756
rect -56 -760 -52 -756
rect -48 -774 -44 -770
rect -40 -774 -36 -770
rect 352 -690 356 -686
rect 360 -690 364 -686
rect 368 -690 372 -686
rect 376 -690 380 -686
rect 289 -704 293 -700
rect 299 -704 303 -700
rect 309 -704 313 -700
rect 324 -704 328 -700
rect 334 -704 338 -700
rect 344 -704 348 -700
rect 253 -718 257 -714
rect 261 -718 265 -714
rect 223 -736 227 -732
rect 231 -736 235 -732
rect 263 -736 267 -732
rect 271 -736 275 -732
rect 279 -736 283 -732
rect 287 -736 291 -732
rect 81 -789 85 -785
rect 91 -789 95 -785
rect 103 -789 107 -785
rect 115 -789 119 -785
rect 125 -789 129 -785
rect -13 -816 -9 -812
rect -5 -816 -1 -812
rect 27 -816 31 -812
rect 35 -816 39 -812
rect 43 -816 47 -812
rect 51 -816 55 -812
rect 151 -853 155 -849
rect 161 -853 165 -849
rect 173 -853 177 -849
rect 185 -853 189 -849
rect 195 -853 199 -849
rect -48 -894 -44 -890
rect -40 -894 -36 -890
rect 15 -886 19 -882
rect 25 -886 29 -882
rect 87 -893 91 -889
rect 98 -893 102 -889
rect 108 -893 112 -889
rect 119 -893 123 -889
rect -13 -903 -9 -899
rect -3 -903 1 -899
rect 7 -903 11 -899
rect -111 -908 -107 -904
rect -101 -908 -97 -904
rect -91 -908 -87 -904
rect -76 -908 -72 -904
rect -66 -908 -62 -904
rect -56 -908 -52 -904
rect -147 -922 -143 -918
rect -139 -922 -135 -918
rect -111 -936 -107 -932
rect -101 -936 -97 -932
rect -91 -936 -87 -932
rect -76 -936 -72 -932
rect -66 -936 -62 -932
rect -56 -936 -52 -932
rect -48 -950 -44 -946
rect -40 -950 -36 -946
rect 87 -980 91 -976
rect 97 -980 101 -976
rect 107 -980 111 -976
rect -147 -1127 -143 -1123
rect -139 -1127 -135 -1123
rect -111 -1141 -107 -1137
rect -101 -1141 -97 -1137
rect -91 -1141 -87 -1137
rect -76 -1141 -72 -1137
rect -66 -1141 -62 -1137
rect -56 -1141 -52 -1137
rect -48 -1155 -44 -1151
rect -40 -1155 -36 -1151
rect 75 -1126 79 -1122
rect 85 -1126 89 -1122
rect 97 -1126 101 -1122
rect 109 -1126 113 -1122
rect 121 -1126 125 -1122
rect 131 -1126 135 -1122
rect -13 -1197 -9 -1193
rect -5 -1197 -1 -1193
rect 27 -1197 31 -1193
rect 35 -1197 39 -1193
rect 43 -1197 47 -1193
rect 51 -1197 55 -1193
rect 321 -1184 325 -1180
rect 329 -1184 333 -1180
rect 337 -1184 341 -1180
rect 345 -1184 349 -1180
rect 258 -1198 262 -1194
rect 268 -1198 272 -1194
rect 293 -1198 297 -1194
rect 303 -1198 307 -1194
rect 313 -1198 317 -1194
rect 83 -1249 87 -1245
rect 93 -1249 97 -1245
rect 105 -1249 109 -1245
rect 117 -1249 121 -1245
rect 127 -1249 131 -1245
rect -48 -1275 -44 -1271
rect -40 -1275 -36 -1271
rect 222 -1212 226 -1208
rect 230 -1212 234 -1208
rect 15 -1267 19 -1263
rect 25 -1267 29 -1263
rect 154 -1266 158 -1262
rect 164 -1266 168 -1262
rect 176 -1266 180 -1262
rect 188 -1266 192 -1262
rect 200 -1266 204 -1262
rect 210 -1266 214 -1262
rect -13 -1284 -9 -1280
rect -3 -1284 1 -1280
rect 7 -1284 11 -1280
rect -111 -1289 -107 -1285
rect -101 -1289 -97 -1285
rect -91 -1289 -87 -1285
rect -76 -1289 -72 -1285
rect -66 -1289 -62 -1285
rect -56 -1289 -52 -1285
rect -147 -1303 -143 -1299
rect -139 -1303 -135 -1299
rect 93 -1355 97 -1351
rect 104 -1355 108 -1351
rect 114 -1355 118 -1351
rect 125 -1355 129 -1351
rect 103 -1443 107 -1439
rect 113 -1443 117 -1439
rect 123 -1443 127 -1439
<< nsubstratencontact >>
rect 55 16 59 20
rect 65 16 69 20
rect 75 16 79 20
rect 91 16 95 20
rect 99 16 103 20
rect 126 16 130 20
rect 134 16 138 20
rect 154 16 158 20
rect 162 16 166 20
rect -20 7 -16 11
rect -12 7 -8 11
rect 252 -8 256 -4
rect 268 -8 272 -4
rect -13 -131 -9 -127
rect -3 -131 1 -127
rect 7 -131 11 -127
rect 58 -131 62 -127
rect 69 -131 73 -127
rect 80 -131 84 -127
rect 90 -131 94 -127
rect 132 -131 136 -127
rect 143 -131 147 -127
rect 154 -131 158 -127
rect 165 -131 169 -127
rect 176 -131 180 -127
rect 240 -131 244 -127
rect 251 -131 255 -127
rect 262 -131 266 -127
rect 273 -131 277 -127
rect 286 -131 290 -127
rect 296 -131 300 -127
rect 27 -331 31 -327
rect 43 -331 47 -327
rect 66 -331 70 -327
rect 76 -331 80 -327
rect 86 -331 90 -327
rect 101 -331 105 -327
rect 111 -331 115 -327
rect 121 -331 125 -327
rect -13 -401 -9 -397
rect -3 -401 1 -397
rect 7 -401 11 -397
rect 15 -401 19 -397
rect 25 -401 29 -397
rect 190 -388 194 -384
rect 206 -388 210 -384
rect -147 -421 -143 -417
rect -137 -421 -133 -417
rect -127 -421 -123 -417
rect -111 -421 -107 -417
rect -103 -421 -99 -417
rect -76 -421 -72 -417
rect -68 -421 -64 -417
rect -48 -421 -44 -417
rect -40 -421 -36 -417
rect 255 -416 259 -412
rect 265 -416 269 -412
rect 275 -416 279 -412
rect 291 -416 295 -412
rect 299 -416 303 -412
rect 326 -416 330 -412
rect 334 -416 338 -412
rect 354 -416 358 -412
rect 362 -416 366 -412
rect 370 -416 374 -412
rect 378 -416 382 -412
rect 75 -478 79 -474
rect 86 -478 90 -474
rect 97 -478 101 -474
rect 107 -478 111 -474
rect 129 -478 133 -474
rect 140 -478 144 -474
rect 151 -478 155 -474
rect 161 -478 165 -474
rect 209 -483 213 -479
rect 225 -483 229 -479
rect 27 -520 31 -516
rect 43 -520 47 -516
rect 75 -582 79 -578
rect 85 -582 89 -578
rect 95 -582 99 -578
rect -13 -590 -9 -586
rect -3 -590 1 -586
rect 7 -590 11 -586
rect 15 -590 19 -586
rect 23 -590 27 -586
rect -147 -597 -143 -593
rect -137 -597 -133 -593
rect -127 -597 -123 -593
rect -111 -597 -107 -593
rect -103 -597 -99 -593
rect -76 -597 -72 -593
rect -68 -597 -64 -593
rect -48 -597 -44 -593
rect -40 -597 -36 -593
rect 253 -630 257 -626
rect 263 -630 267 -626
rect 273 -630 277 -626
rect 289 -630 293 -626
rect 297 -630 301 -626
rect 324 -630 328 -626
rect 332 -630 336 -626
rect 352 -630 356 -626
rect 360 -630 364 -626
rect 368 -630 372 -626
rect 376 -630 380 -626
rect 81 -678 85 -674
rect 92 -678 96 -674
rect 103 -678 107 -674
rect 114 -678 118 -674
rect 125 -678 129 -674
rect 191 -710 195 -706
rect 207 -710 211 -706
rect 27 -756 31 -752
rect 43 -756 47 -752
rect 151 -742 155 -738
rect 162 -742 166 -738
rect 173 -742 177 -738
rect 184 -742 188 -738
rect 195 -742 199 -738
rect 87 -799 91 -795
rect 98 -799 102 -795
rect 109 -799 113 -795
rect 119 -799 123 -795
rect -13 -826 -9 -822
rect -3 -826 1 -822
rect 7 -826 11 -822
rect 15 -826 19 -822
rect 25 -826 29 -822
rect -147 -834 -143 -830
rect -137 -834 -133 -830
rect -127 -834 -123 -830
rect -111 -834 -107 -830
rect -103 -834 -99 -830
rect -76 -834 -72 -830
rect -68 -834 -64 -830
rect -48 -834 -44 -830
rect -40 -834 -36 -830
rect 263 -796 267 -792
rect 279 -796 283 -792
rect 87 -903 91 -899
rect 97 -903 101 -899
rect 107 -903 111 -899
rect 75 -998 79 -994
rect 86 -998 90 -994
rect 97 -998 101 -994
rect 108 -998 112 -994
rect 121 -998 125 -994
rect 131 -998 135 -994
rect -147 -1010 -143 -1006
rect -137 -1010 -133 -1006
rect -127 -1010 -123 -1006
rect -111 -1010 -107 -1006
rect -103 -1010 -99 -1006
rect -76 -1010 -72 -1006
rect -68 -1010 -64 -1006
rect -48 -1010 -44 -1006
rect -40 -1010 -36 -1006
rect 222 -1124 226 -1120
rect 232 -1124 236 -1120
rect 242 -1124 246 -1120
rect 258 -1124 262 -1120
rect 266 -1124 270 -1120
rect 293 -1124 297 -1120
rect 301 -1124 305 -1120
rect 321 -1124 325 -1120
rect 329 -1124 333 -1120
rect 337 -1124 341 -1120
rect 345 -1124 349 -1120
rect 27 -1137 31 -1133
rect 43 -1137 47 -1133
rect 83 -1138 87 -1134
rect 94 -1138 98 -1134
rect 105 -1138 109 -1134
rect 116 -1138 120 -1134
rect 127 -1138 131 -1134
rect 154 -1138 158 -1134
rect 165 -1138 169 -1134
rect 176 -1138 180 -1134
rect 187 -1138 191 -1134
rect 200 -1138 204 -1134
rect 210 -1138 214 -1134
rect -13 -1207 -9 -1203
rect -3 -1207 1 -1203
rect 7 -1207 11 -1203
rect 15 -1207 19 -1203
rect 25 -1207 29 -1203
rect -147 -1215 -143 -1211
rect -137 -1215 -133 -1211
rect -127 -1215 -123 -1211
rect -111 -1215 -107 -1211
rect -103 -1215 -99 -1211
rect -76 -1215 -72 -1211
rect -68 -1215 -64 -1211
rect -48 -1215 -44 -1211
rect -40 -1215 -36 -1211
rect 93 -1261 97 -1257
rect 104 -1261 108 -1257
rect 115 -1261 119 -1257
rect 125 -1261 129 -1257
rect 103 -1366 107 -1362
rect 113 -1366 117 -1362
rect 123 -1366 127 -1362
<< polysilicon >>
rect 60 10 62 13
rect 72 10 74 13
rect 96 10 98 13
rect 131 10 133 13
rect 159 10 161 13
rect 217 11 219 14
rect 233 11 235 14
rect -15 1 -13 4
rect -15 -35 -13 -19
rect 96 -30 98 -10
rect 108 -30 110 -23
rect 131 -30 133 -10
rect 143 -30 145 -23
rect 159 -26 161 -10
rect -15 -48 -13 -45
rect 60 -54 62 -30
rect 72 -44 74 -30
rect 257 -14 259 -11
rect 273 -14 275 -11
rect 159 -39 161 -36
rect 217 -50 219 -29
rect 233 -40 235 -29
rect 257 -50 259 -34
rect 273 -50 275 -34
rect 96 -53 98 -50
rect 108 -53 110 -50
rect 131 -53 133 -50
rect 143 -53 145 -50
rect 217 -63 219 -60
rect 257 -63 259 -60
rect 273 -63 275 -60
rect 60 -67 62 -64
rect -8 -137 -6 -134
rect 4 -137 6 -134
rect 63 -137 65 -134
rect 75 -137 77 -134
rect 87 -137 89 -134
rect 137 -137 139 -134
rect 149 -137 151 -134
rect 161 -137 163 -134
rect 173 -137 175 -134
rect 245 -137 247 -134
rect 257 -137 259 -134
rect 269 -137 271 -134
rect 281 -137 283 -134
rect 293 -137 295 -134
rect -8 -180 -6 -157
rect 4 -180 6 -157
rect 63 -187 65 -157
rect 75 -187 77 -157
rect 87 -187 89 -157
rect -8 -203 -6 -200
rect 4 -203 6 -200
rect 137 -194 139 -157
rect 149 -194 151 -157
rect 161 -194 163 -157
rect 173 -194 175 -157
rect 63 -220 65 -217
rect 75 -220 77 -217
rect 87 -220 89 -217
rect 245 -201 247 -157
rect 257 -201 259 -157
rect 269 -201 271 -157
rect 281 -201 283 -157
rect 293 -201 295 -157
rect 137 -237 139 -234
rect 149 -237 151 -234
rect 161 -237 163 -234
rect 173 -237 175 -234
rect 245 -254 247 -251
rect 257 -254 259 -251
rect 269 -254 271 -251
rect 281 -254 283 -251
rect 293 -254 295 -251
rect -8 -312 -6 -309
rect 8 -312 10 -309
rect -142 -337 -140 -334
rect -142 -371 -140 -347
rect -106 -351 -104 -348
rect -94 -351 -92 -348
rect -71 -351 -69 -348
rect -59 -351 -57 -348
rect -130 -371 -128 -357
rect 155 -332 157 -329
rect 195 -332 197 -329
rect 211 -332 213 -329
rect 260 -332 262 -329
rect 32 -337 34 -334
rect 48 -337 50 -334
rect 71 -337 73 -334
rect 83 -337 85 -334
rect 106 -337 108 -334
rect 118 -337 120 -334
rect -43 -365 -41 -362
rect -106 -391 -104 -371
rect -94 -378 -92 -371
rect -71 -391 -69 -371
rect -59 -378 -57 -371
rect -8 -373 -6 -352
rect 8 -363 10 -352
rect 32 -373 34 -357
rect 48 -373 50 -357
rect -43 -391 -41 -375
rect 71 -380 73 -357
rect 83 -380 85 -357
rect 106 -380 108 -357
rect 118 -380 120 -357
rect 155 -363 157 -342
rect 171 -363 173 -352
rect 195 -358 197 -342
rect 211 -358 213 -342
rect -8 -386 -6 -383
rect 32 -386 34 -383
rect 48 -386 50 -383
rect 71 -403 73 -400
rect 83 -403 85 -400
rect 106 -403 108 -400
rect 118 -403 120 -400
rect 260 -366 262 -342
rect 296 -346 298 -343
rect 308 -346 310 -343
rect 331 -346 333 -343
rect 343 -346 345 -343
rect 272 -366 274 -352
rect 359 -360 361 -357
rect 375 -360 377 -357
rect 195 -381 197 -378
rect 211 -381 213 -378
rect -8 -407 -6 -404
rect 4 -407 6 -404
rect 20 -407 22 -404
rect -142 -414 -140 -411
rect -130 -414 -128 -411
rect -106 -414 -104 -411
rect -71 -414 -69 -411
rect -43 -414 -41 -411
rect -142 -427 -140 -424
rect -130 -427 -128 -424
rect -106 -427 -104 -424
rect -71 -427 -69 -424
rect -43 -427 -41 -424
rect 155 -406 157 -403
rect 171 -406 173 -403
rect 296 -386 298 -366
rect 308 -373 310 -366
rect 331 -386 333 -366
rect 343 -373 345 -366
rect 359 -386 361 -370
rect 375 -386 377 -370
rect 260 -409 262 -406
rect 272 -409 274 -406
rect 296 -409 298 -406
rect 331 -409 333 -406
rect 359 -409 361 -406
rect 375 -409 377 -406
rect 260 -422 262 -419
rect 272 -422 274 -419
rect 296 -422 298 -419
rect 331 -422 333 -419
rect 359 -422 361 -419
rect 375 -422 377 -419
rect 174 -427 176 -424
rect 214 -427 216 -424
rect 230 -427 232 -424
rect -106 -467 -104 -447
rect -94 -467 -92 -460
rect -71 -467 -69 -447
rect -59 -467 -57 -460
rect -43 -463 -41 -447
rect -8 -450 -6 -427
rect 4 -450 6 -427
rect 20 -443 22 -427
rect -142 -491 -140 -467
rect -130 -481 -128 -467
rect 20 -456 22 -453
rect 174 -458 176 -437
rect 190 -458 192 -447
rect 214 -453 216 -437
rect 230 -453 232 -437
rect -8 -473 -6 -470
rect 4 -473 6 -470
rect -43 -476 -41 -473
rect 80 -484 82 -481
rect 92 -484 94 -481
rect 104 -484 106 -481
rect 134 -484 136 -481
rect 146 -484 148 -481
rect 158 -484 160 -481
rect -106 -490 -104 -487
rect -94 -490 -92 -487
rect -71 -490 -69 -487
rect -59 -490 -57 -487
rect -8 -501 -6 -498
rect 8 -501 10 -498
rect -142 -504 -140 -501
rect -142 -513 -140 -510
rect -142 -547 -140 -523
rect -106 -527 -104 -524
rect -94 -527 -92 -524
rect -71 -527 -69 -524
rect -59 -527 -57 -524
rect -130 -547 -128 -533
rect -43 -541 -41 -538
rect 296 -462 298 -442
rect 308 -462 310 -455
rect 331 -462 333 -442
rect 343 -462 345 -455
rect 359 -458 361 -442
rect 375 -458 377 -442
rect 214 -476 216 -473
rect 230 -476 232 -473
rect 260 -486 262 -462
rect 272 -476 274 -462
rect 359 -471 361 -468
rect 375 -471 377 -468
rect 296 -485 298 -482
rect 308 -485 310 -482
rect 331 -485 333 -482
rect 343 -485 345 -482
rect 174 -501 176 -498
rect 190 -501 192 -498
rect 260 -499 262 -496
rect 32 -526 34 -523
rect 48 -526 50 -523
rect -106 -567 -104 -547
rect -94 -554 -92 -547
rect -71 -567 -69 -547
rect -59 -554 -57 -547
rect -43 -567 -41 -551
rect -8 -562 -6 -541
rect 8 -552 10 -541
rect 80 -534 82 -504
rect 92 -534 94 -504
rect 104 -534 106 -504
rect 134 -534 136 -504
rect 146 -534 148 -504
rect 158 -534 160 -504
rect 32 -562 34 -546
rect 48 -562 50 -546
rect 258 -546 260 -543
rect 80 -567 82 -564
rect 92 -567 94 -564
rect 104 -567 106 -564
rect 134 -567 136 -564
rect 146 -567 148 -564
rect 158 -567 160 -564
rect -8 -575 -6 -572
rect 32 -575 34 -572
rect 48 -575 50 -572
rect 258 -580 260 -556
rect 294 -560 296 -557
rect 306 -560 308 -557
rect 329 -560 331 -557
rect 341 -560 343 -557
rect 270 -580 272 -566
rect 357 -574 359 -571
rect 373 -574 375 -571
rect -142 -590 -140 -587
rect -130 -590 -128 -587
rect -106 -590 -104 -587
rect -71 -590 -69 -587
rect -43 -590 -41 -587
rect 80 -588 82 -585
rect 92 -588 94 -585
rect -8 -596 -6 -593
rect 4 -596 6 -593
rect 20 -596 22 -593
rect -142 -603 -140 -600
rect -130 -603 -128 -600
rect -106 -603 -104 -600
rect -71 -603 -69 -600
rect -43 -603 -41 -600
rect -106 -643 -104 -623
rect -94 -643 -92 -636
rect -71 -643 -69 -623
rect -59 -643 -57 -636
rect -43 -639 -41 -623
rect -8 -639 -6 -616
rect 4 -639 6 -616
rect 20 -632 22 -616
rect 80 -631 82 -608
rect 92 -631 94 -608
rect 294 -600 296 -580
rect 306 -587 308 -580
rect 329 -600 331 -580
rect 341 -587 343 -580
rect 357 -600 359 -584
rect 373 -600 375 -584
rect 258 -623 260 -620
rect 270 -623 272 -620
rect 294 -623 296 -620
rect 329 -623 331 -620
rect 357 -623 359 -620
rect 373 -623 375 -620
rect -142 -667 -140 -643
rect -130 -657 -128 -643
rect -43 -652 -41 -649
rect 20 -645 22 -642
rect 258 -636 260 -633
rect 270 -636 272 -633
rect 294 -636 296 -633
rect 329 -636 331 -633
rect 357 -636 359 -633
rect 373 -636 375 -633
rect 80 -654 82 -651
rect 92 -654 94 -651
rect 156 -654 158 -651
rect 196 -654 198 -651
rect 212 -654 214 -651
rect -8 -662 -6 -659
rect 4 -662 6 -659
rect -106 -666 -104 -663
rect -94 -666 -92 -663
rect -71 -666 -69 -663
rect -59 -666 -57 -663
rect -142 -680 -140 -677
rect 86 -684 88 -681
rect 98 -684 100 -681
rect 110 -684 112 -681
rect 122 -684 124 -681
rect 156 -685 158 -664
rect 172 -685 174 -674
rect 196 -680 198 -664
rect 212 -680 214 -664
rect 294 -676 296 -656
rect 306 -676 308 -669
rect 329 -676 331 -656
rect 341 -676 343 -669
rect 357 -672 359 -656
rect 373 -672 375 -656
rect -8 -737 -6 -734
rect 8 -737 10 -734
rect -142 -750 -140 -747
rect -142 -784 -140 -760
rect -106 -764 -104 -761
rect -94 -764 -92 -761
rect -71 -764 -69 -761
rect -59 -764 -57 -761
rect -130 -784 -128 -770
rect -43 -778 -41 -775
rect 86 -741 88 -704
rect 98 -741 100 -704
rect 110 -741 112 -704
rect 122 -741 124 -704
rect 258 -700 260 -676
rect 270 -690 272 -676
rect 357 -685 359 -682
rect 373 -685 375 -682
rect 294 -699 296 -696
rect 306 -699 308 -696
rect 329 -699 331 -696
rect 341 -699 343 -696
rect 196 -703 198 -700
rect 212 -703 214 -700
rect 258 -713 260 -710
rect 156 -728 158 -725
rect 172 -728 174 -725
rect 32 -762 34 -759
rect 48 -762 50 -759
rect -106 -804 -104 -784
rect -94 -791 -92 -784
rect -71 -804 -69 -784
rect -59 -791 -57 -784
rect -43 -804 -41 -788
rect -8 -798 -6 -777
rect 8 -788 10 -777
rect 228 -740 230 -737
rect 268 -740 270 -737
rect 284 -740 286 -737
rect 156 -748 158 -745
rect 168 -748 170 -745
rect 180 -748 182 -745
rect 192 -748 194 -745
rect 32 -798 34 -782
rect 48 -798 50 -782
rect 86 -784 88 -781
rect 98 -784 100 -781
rect 110 -784 112 -781
rect 122 -784 124 -781
rect 92 -805 94 -802
rect 104 -805 106 -802
rect 116 -805 118 -802
rect 156 -805 158 -768
rect 168 -805 170 -768
rect 180 -805 182 -768
rect 192 -805 194 -768
rect 228 -771 230 -750
rect 244 -771 246 -760
rect 268 -766 270 -750
rect 284 -766 286 -750
rect -8 -811 -6 -808
rect 32 -811 34 -808
rect 48 -811 50 -808
rect -142 -827 -140 -824
rect -130 -827 -128 -824
rect -106 -827 -104 -824
rect -71 -827 -69 -824
rect -43 -827 -41 -824
rect -8 -832 -6 -829
rect 4 -832 6 -829
rect 20 -832 22 -829
rect -142 -840 -140 -837
rect -130 -840 -128 -837
rect -106 -840 -104 -837
rect -71 -840 -69 -837
rect -43 -840 -41 -837
rect -106 -880 -104 -860
rect -94 -880 -92 -873
rect -71 -880 -69 -860
rect -59 -880 -57 -873
rect -43 -876 -41 -860
rect -8 -875 -6 -852
rect 4 -875 6 -852
rect 20 -868 22 -852
rect 92 -855 94 -825
rect 104 -855 106 -825
rect 116 -855 118 -825
rect 268 -789 270 -786
rect 284 -789 286 -786
rect 228 -814 230 -811
rect 244 -814 246 -811
rect 156 -848 158 -845
rect 168 -848 170 -845
rect 180 -848 182 -845
rect 192 -848 194 -845
rect -142 -904 -140 -880
rect -130 -894 -128 -880
rect -43 -889 -41 -886
rect 20 -881 22 -878
rect 92 -888 94 -885
rect 104 -888 106 -885
rect 116 -888 118 -885
rect -8 -898 -6 -895
rect 4 -898 6 -895
rect -106 -903 -104 -900
rect -94 -903 -92 -900
rect -71 -903 -69 -900
rect -59 -903 -57 -900
rect 92 -909 94 -906
rect 104 -909 106 -906
rect -142 -917 -140 -914
rect -142 -926 -140 -923
rect -142 -960 -140 -936
rect -106 -940 -104 -937
rect -94 -940 -92 -937
rect -71 -940 -69 -937
rect -59 -940 -57 -937
rect -130 -960 -128 -946
rect -43 -954 -41 -951
rect 92 -952 94 -929
rect 104 -952 106 -929
rect -106 -980 -104 -960
rect -94 -967 -92 -960
rect -71 -980 -69 -960
rect -59 -967 -57 -960
rect -43 -980 -41 -964
rect 92 -975 94 -972
rect 104 -975 106 -972
rect -142 -1003 -140 -1000
rect -130 -1003 -128 -1000
rect -106 -1003 -104 -1000
rect -71 -1003 -69 -1000
rect -43 -1003 -41 -1000
rect 80 -1004 82 -1001
rect 92 -1004 94 -1001
rect 104 -1004 106 -1001
rect 116 -1004 118 -1001
rect 128 -1004 130 -1001
rect 80 -1068 82 -1024
rect 92 -1068 94 -1024
rect 104 -1068 106 -1024
rect 116 -1068 118 -1024
rect 128 -1068 130 -1024
rect -8 -1118 -6 -1115
rect 8 -1118 10 -1115
rect -142 -1131 -140 -1128
rect -142 -1165 -140 -1141
rect -106 -1145 -104 -1142
rect -94 -1145 -92 -1142
rect -71 -1145 -69 -1142
rect -59 -1145 -57 -1142
rect -130 -1165 -128 -1151
rect -43 -1159 -41 -1156
rect 80 -1121 82 -1118
rect 92 -1121 94 -1118
rect 104 -1121 106 -1118
rect 116 -1121 118 -1118
rect 128 -1121 130 -1118
rect 227 -1130 229 -1127
rect 239 -1130 241 -1127
rect 263 -1130 265 -1127
rect 298 -1130 300 -1127
rect 326 -1130 328 -1127
rect 342 -1130 344 -1127
rect 32 -1143 34 -1140
rect 48 -1143 50 -1140
rect -106 -1185 -104 -1165
rect -94 -1172 -92 -1165
rect -71 -1185 -69 -1165
rect -59 -1172 -57 -1165
rect -43 -1185 -41 -1169
rect -8 -1179 -6 -1158
rect 8 -1169 10 -1158
rect 88 -1144 90 -1141
rect 100 -1144 102 -1141
rect 112 -1144 114 -1141
rect 124 -1144 126 -1141
rect 159 -1144 161 -1141
rect 171 -1144 173 -1141
rect 183 -1144 185 -1141
rect 195 -1144 197 -1141
rect 207 -1144 209 -1141
rect 32 -1179 34 -1163
rect 48 -1179 50 -1163
rect -8 -1192 -6 -1189
rect 32 -1192 34 -1189
rect 48 -1192 50 -1189
rect 88 -1201 90 -1164
rect 100 -1201 102 -1164
rect 112 -1201 114 -1164
rect 124 -1201 126 -1164
rect -142 -1208 -140 -1205
rect -130 -1208 -128 -1205
rect -106 -1208 -104 -1205
rect -71 -1208 -69 -1205
rect -43 -1208 -41 -1205
rect -8 -1213 -6 -1210
rect 4 -1213 6 -1210
rect 20 -1213 22 -1210
rect -142 -1221 -140 -1218
rect -130 -1221 -128 -1218
rect -106 -1221 -104 -1218
rect -71 -1221 -69 -1218
rect -43 -1221 -41 -1218
rect -106 -1261 -104 -1241
rect -94 -1261 -92 -1254
rect -71 -1261 -69 -1241
rect -59 -1261 -57 -1254
rect -43 -1257 -41 -1241
rect -8 -1256 -6 -1233
rect 4 -1256 6 -1233
rect 20 -1249 22 -1233
rect 159 -1208 161 -1164
rect 171 -1208 173 -1164
rect 183 -1208 185 -1164
rect 195 -1208 197 -1164
rect 207 -1208 209 -1164
rect 263 -1170 265 -1150
rect 275 -1170 277 -1163
rect 298 -1170 300 -1150
rect 310 -1170 312 -1163
rect 326 -1166 328 -1150
rect 342 -1166 344 -1150
rect 227 -1194 229 -1170
rect 239 -1184 241 -1170
rect 326 -1179 328 -1176
rect 342 -1179 344 -1176
rect 263 -1193 265 -1190
rect 275 -1193 277 -1190
rect 298 -1193 300 -1190
rect 310 -1193 312 -1190
rect 227 -1207 229 -1204
rect 88 -1244 90 -1241
rect 100 -1244 102 -1241
rect 112 -1244 114 -1241
rect 124 -1244 126 -1241
rect -142 -1285 -140 -1261
rect -130 -1275 -128 -1261
rect -43 -1270 -41 -1267
rect 20 -1262 22 -1259
rect 159 -1261 161 -1258
rect 171 -1261 173 -1258
rect 183 -1261 185 -1258
rect 195 -1261 197 -1258
rect 207 -1261 209 -1258
rect 98 -1267 100 -1264
rect 110 -1267 112 -1264
rect 122 -1267 124 -1264
rect -8 -1279 -6 -1276
rect 4 -1279 6 -1276
rect -106 -1284 -104 -1281
rect -94 -1284 -92 -1281
rect -71 -1284 -69 -1281
rect -59 -1284 -57 -1281
rect -142 -1298 -140 -1295
rect 98 -1317 100 -1287
rect 110 -1317 112 -1287
rect 122 -1317 124 -1287
rect 98 -1350 100 -1347
rect 110 -1350 112 -1347
rect 122 -1350 124 -1347
rect 108 -1372 110 -1369
rect 120 -1372 122 -1369
rect 108 -1415 110 -1392
rect 120 -1415 122 -1392
rect 108 -1438 110 -1435
rect 120 -1438 122 -1435
<< polycontact >>
rect -19 -32 -15 -28
rect 92 -20 96 -16
rect 127 -21 131 -17
rect 104 -27 108 -23
rect 155 -23 159 -19
rect 139 -27 143 -23
rect 56 -51 60 -47
rect 68 -42 72 -38
rect 213 -47 217 -43
rect 229 -40 233 -36
rect 253 -47 257 -43
rect 269 -47 273 -43
rect -12 -170 -8 -166
rect 0 -177 4 -173
rect 59 -170 63 -166
rect 71 -177 75 -173
rect 83 -184 87 -180
rect 133 -170 137 -166
rect 145 -177 149 -173
rect 157 -184 161 -180
rect 169 -191 173 -187
rect 241 -170 245 -166
rect 253 -177 257 -173
rect 265 -184 269 -180
rect 277 -191 281 -187
rect 289 -198 293 -194
rect -146 -354 -142 -350
rect -134 -363 -130 -359
rect -110 -385 -106 -381
rect -98 -378 -94 -374
rect -75 -384 -71 -380
rect -63 -378 -59 -374
rect -12 -370 -8 -366
rect 4 -363 8 -359
rect 151 -349 155 -345
rect 28 -370 32 -366
rect 44 -370 48 -366
rect 67 -370 71 -366
rect -47 -382 -43 -378
rect 79 -377 83 -373
rect 102 -370 106 -366
rect 114 -377 118 -373
rect 191 -349 195 -345
rect 167 -356 171 -352
rect 207 -349 211 -345
rect 256 -349 260 -345
rect 268 -358 272 -354
rect 292 -380 296 -376
rect 304 -373 308 -369
rect 327 -379 331 -375
rect 339 -373 343 -369
rect 355 -377 359 -373
rect 371 -377 375 -373
rect -12 -440 -8 -436
rect -110 -457 -106 -453
rect -75 -458 -71 -454
rect -98 -464 -94 -460
rect -47 -460 -43 -456
rect -63 -464 -59 -460
rect 0 -447 4 -443
rect 16 -440 20 -436
rect -146 -488 -142 -484
rect -134 -479 -130 -475
rect 170 -444 174 -440
rect 210 -444 214 -440
rect 186 -451 190 -447
rect 226 -444 230 -440
rect -146 -530 -142 -526
rect -134 -539 -130 -535
rect 292 -452 296 -448
rect 327 -453 331 -449
rect 304 -459 308 -455
rect 355 -455 359 -451
rect 339 -459 343 -455
rect 371 -455 375 -451
rect 256 -483 260 -479
rect 268 -474 272 -470
rect 76 -517 80 -513
rect -110 -561 -106 -557
rect -98 -554 -94 -550
rect -75 -560 -71 -556
rect -63 -554 -59 -550
rect -47 -558 -43 -554
rect -12 -559 -8 -555
rect 4 -552 8 -548
rect 88 -524 92 -520
rect 100 -531 104 -527
rect 130 -517 134 -513
rect 142 -524 146 -520
rect 154 -531 158 -527
rect 28 -559 32 -555
rect 44 -559 48 -555
rect 254 -563 258 -559
rect 266 -572 270 -568
rect -110 -633 -106 -629
rect -75 -634 -71 -630
rect -98 -640 -94 -636
rect -47 -636 -43 -632
rect -63 -640 -59 -636
rect -12 -629 -8 -625
rect 0 -636 4 -632
rect 16 -629 20 -625
rect 76 -621 80 -617
rect 88 -628 92 -624
rect 290 -594 294 -590
rect 302 -587 306 -583
rect 325 -593 329 -589
rect 337 -587 341 -583
rect 353 -591 357 -587
rect 369 -591 373 -587
rect -146 -664 -142 -660
rect -134 -655 -130 -651
rect 152 -671 156 -667
rect 192 -671 196 -667
rect 168 -678 172 -674
rect 208 -671 212 -667
rect 290 -666 294 -662
rect 325 -667 329 -663
rect 302 -673 306 -669
rect 353 -669 357 -665
rect 337 -673 341 -669
rect 369 -669 373 -665
rect 82 -717 86 -713
rect -146 -767 -142 -763
rect -134 -776 -130 -772
rect 94 -724 98 -720
rect 106 -731 110 -727
rect 118 -738 122 -734
rect 254 -697 258 -693
rect 266 -688 270 -684
rect -110 -798 -106 -794
rect -98 -791 -94 -787
rect -75 -797 -71 -793
rect -63 -791 -59 -787
rect -47 -795 -43 -791
rect -12 -795 -8 -791
rect 4 -788 8 -784
rect 224 -757 228 -753
rect 152 -781 156 -777
rect 28 -795 32 -791
rect 44 -795 48 -791
rect 164 -788 168 -784
rect 176 -795 180 -791
rect 188 -802 192 -798
rect 264 -757 268 -753
rect 240 -764 244 -760
rect 280 -757 284 -753
rect 88 -838 92 -834
rect -110 -870 -106 -866
rect -75 -871 -71 -867
rect -98 -877 -94 -873
rect -47 -873 -43 -869
rect -63 -877 -59 -873
rect -12 -865 -8 -861
rect 0 -872 4 -868
rect 16 -865 20 -861
rect 100 -845 104 -841
rect 112 -852 116 -848
rect -146 -901 -142 -897
rect -134 -892 -130 -888
rect -146 -943 -142 -939
rect -134 -952 -130 -948
rect 88 -942 92 -938
rect 100 -949 104 -945
rect -110 -974 -106 -970
rect -98 -967 -94 -963
rect -75 -973 -71 -969
rect -63 -967 -59 -963
rect -47 -971 -43 -967
rect 76 -1037 80 -1033
rect 88 -1044 92 -1040
rect 100 -1051 104 -1047
rect 112 -1058 116 -1054
rect 124 -1065 128 -1061
rect -146 -1148 -142 -1144
rect -134 -1157 -130 -1153
rect -110 -1179 -106 -1175
rect -98 -1172 -94 -1168
rect -75 -1178 -71 -1174
rect -63 -1172 -59 -1168
rect -47 -1176 -43 -1172
rect -12 -1176 -8 -1172
rect 4 -1169 8 -1165
rect 28 -1176 32 -1172
rect 44 -1176 48 -1172
rect 84 -1177 88 -1173
rect 96 -1184 100 -1180
rect 108 -1191 112 -1187
rect 120 -1198 124 -1194
rect 155 -1177 159 -1173
rect -110 -1251 -106 -1247
rect -75 -1252 -71 -1248
rect -98 -1258 -94 -1254
rect -47 -1254 -43 -1250
rect -63 -1258 -59 -1254
rect -12 -1246 -8 -1242
rect 0 -1253 4 -1249
rect 16 -1246 20 -1242
rect 167 -1184 171 -1180
rect 179 -1191 183 -1187
rect 191 -1198 195 -1194
rect 203 -1205 207 -1201
rect 259 -1160 263 -1156
rect 294 -1161 298 -1157
rect 271 -1167 275 -1163
rect 322 -1163 326 -1159
rect 306 -1167 310 -1163
rect 338 -1163 342 -1159
rect 223 -1191 227 -1187
rect 235 -1182 239 -1178
rect -146 -1282 -142 -1278
rect -134 -1273 -130 -1269
rect 94 -1300 98 -1296
rect 106 -1307 110 -1303
rect 118 -1314 122 -1310
rect 104 -1405 108 -1401
rect 116 -1412 120 -1408
<< metal1 >>
rect 59 16 65 20
rect 69 16 75 20
rect 79 16 91 20
rect 95 16 99 20
rect 103 16 126 20
rect 130 16 134 20
rect 138 16 154 20
rect 158 16 162 20
rect 212 17 246 21
rect -16 7 -12 11
rect 55 10 59 16
rect 91 10 95 16
rect 126 10 130 16
rect 154 10 158 16
rect 212 11 216 17
rect 228 11 232 17
rect -20 1 -16 7
rect -12 -28 -8 -19
rect -26 -32 -19 -28
rect -12 -32 -2 -28
rect 90 -20 92 -16
rect 99 -17 103 -10
rect 134 -17 138 -10
rect 99 -20 127 -17
rect 111 -21 127 -20
rect 134 -19 150 -17
rect 162 -19 166 -10
rect 134 -20 155 -19
rect 79 -27 104 -24
rect 111 -30 115 -21
rect 146 -23 155 -20
rect 162 -23 172 -19
rect 123 -27 139 -24
rect 146 -30 150 -23
rect 162 -26 166 -23
rect -12 -35 -8 -32
rect 49 -42 53 -38
rect 58 -42 68 -38
rect -20 -49 -16 -45
rect 75 -47 79 -30
rect -16 -53 -12 -49
rect 49 -51 56 -47
rect 63 -51 79 -47
rect 221 -36 224 -29
rect 154 -40 158 -36
rect 206 -40 229 -36
rect 158 -44 162 -40
rect 237 -43 240 -29
rect 63 -54 67 -51
rect 91 -54 95 -50
rect 126 -54 130 -50
rect 154 -54 158 -44
rect 206 -47 213 -43
rect 217 -47 240 -43
rect 243 -43 246 17
rect 256 -8 268 -4
rect 252 -14 256 -8
rect 268 -14 272 -8
rect 260 -43 264 -34
rect 276 -43 280 -34
rect 243 -47 253 -43
rect 260 -47 269 -43
rect 276 -47 286 -43
rect 243 -50 246 -47
rect 260 -50 264 -47
rect 276 -50 280 -47
rect 72 -58 91 -54
rect 95 -58 101 -54
rect 105 -58 126 -54
rect 130 -58 136 -54
rect 140 -58 146 -54
rect 150 -58 158 -54
rect 55 -68 59 -64
rect 72 -68 76 -58
rect 224 -53 246 -50
rect 212 -64 216 -60
rect 252 -64 256 -60
rect 268 -64 272 -60
rect 216 -68 220 -64
rect 224 -68 252 -64
rect 256 -68 260 -64
rect 264 -68 268 -64
rect 272 -68 276 -64
rect 59 -72 63 -68
rect 67 -72 76 -68
rect -9 -131 -3 -127
rect 1 -131 7 -127
rect -13 -137 -9 -131
rect 7 -137 11 -131
rect 62 -131 69 -127
rect 73 -131 80 -127
rect 84 -131 90 -127
rect 136 -131 143 -127
rect 147 -131 154 -127
rect 158 -131 165 -127
rect 169 -131 176 -127
rect 58 -137 62 -131
rect 80 -137 84 -131
rect 132 -137 136 -131
rect 154 -137 158 -131
rect 176 -137 180 -131
rect 244 -131 251 -127
rect 255 -131 262 -127
rect 266 -131 273 -127
rect 277 -131 286 -127
rect 290 -131 296 -127
rect 240 -137 244 -131
rect 262 -137 266 -131
rect 286 -137 290 -131
rect -3 -166 1 -157
rect 68 -166 72 -157
rect 90 -166 94 -157
rect 142 -160 146 -157
rect 166 -160 170 -157
rect 142 -163 170 -160
rect 250 -160 254 -157
rect 274 -160 278 -157
rect 296 -160 300 -157
rect 250 -163 300 -160
rect -19 -170 -12 -166
rect -3 -170 17 -166
rect 52 -170 59 -166
rect 68 -170 94 -166
rect 126 -170 133 -166
rect -19 -177 0 -173
rect 7 -180 11 -170
rect 90 -173 94 -170
rect 166 -173 170 -163
rect 234 -170 241 -166
rect 52 -177 71 -173
rect 90 -177 100 -173
rect 126 -177 145 -173
rect 166 -177 186 -173
rect 234 -177 253 -173
rect 52 -184 83 -180
rect 90 -187 94 -177
rect 126 -184 157 -180
rect -13 -204 -9 -200
rect -9 -208 -3 -204
rect 1 -208 7 -204
rect 126 -191 169 -187
rect 176 -194 180 -177
rect 296 -180 300 -163
rect 234 -184 265 -180
rect 296 -184 306 -180
rect 234 -191 277 -187
rect 58 -221 62 -217
rect 62 -225 69 -221
rect 73 -225 79 -221
rect 83 -225 90 -221
rect 234 -198 289 -194
rect 296 -201 300 -184
rect 132 -238 136 -234
rect 136 -242 142 -238
rect 146 -242 154 -238
rect 158 -242 166 -238
rect 170 -242 176 -238
rect 240 -255 244 -251
rect 244 -259 250 -255
rect 254 -259 262 -255
rect 266 -259 274 -255
rect 278 -259 286 -255
rect 290 -259 296 -255
rect -13 -306 21 -302
rect -13 -312 -9 -306
rect 3 -312 7 -306
rect -143 -333 -139 -329
rect -135 -333 -126 -329
rect -147 -337 -143 -333
rect -130 -343 -126 -333
rect -130 -347 -111 -343
rect -107 -347 -101 -343
rect -97 -347 -91 -343
rect -87 -347 -76 -343
rect -72 -347 -66 -343
rect -62 -347 -56 -343
rect -52 -347 -44 -343
rect -139 -350 -135 -347
rect -153 -354 -146 -350
rect -139 -354 -123 -350
rect -148 -363 -134 -359
rect -127 -371 -123 -354
rect -111 -351 -107 -347
rect -76 -351 -72 -347
rect -123 -377 -98 -374
rect -91 -380 -87 -371
rect -79 -377 -63 -374
rect -56 -378 -52 -371
rect -48 -357 -44 -347
rect -44 -361 -40 -357
rect -4 -359 -1 -352
rect -48 -365 -44 -361
rect -27 -362 4 -359
rect -40 -378 -36 -375
rect -27 -378 -24 -362
rect 12 -366 15 -352
rect -16 -370 -12 -366
rect -8 -370 15 -366
rect 18 -366 21 -306
rect 31 -331 43 -327
rect 27 -337 31 -331
rect 43 -337 47 -331
rect 70 -331 76 -327
rect 80 -331 86 -327
rect 90 -330 101 -327
rect 66 -337 70 -331
rect 86 -337 90 -331
rect 105 -331 111 -327
rect 115 -331 121 -327
rect 101 -337 105 -331
rect 121 -337 125 -331
rect 154 -328 158 -324
rect 162 -328 190 -324
rect 194 -328 198 -324
rect 202 -328 206 -324
rect 210 -328 214 -324
rect 259 -328 263 -324
rect 267 -328 276 -324
rect 150 -332 154 -328
rect 190 -332 194 -328
rect 206 -332 210 -328
rect 255 -332 259 -328
rect 162 -342 184 -339
rect 272 -338 276 -328
rect 272 -342 291 -338
rect 295 -342 301 -338
rect 305 -342 311 -338
rect 315 -342 326 -338
rect 330 -342 336 -338
rect 340 -342 346 -338
rect 350 -342 358 -338
rect 181 -345 184 -342
rect 198 -345 202 -342
rect 214 -345 218 -342
rect 263 -345 267 -342
rect 137 -349 151 -345
rect 155 -349 178 -345
rect 144 -356 167 -352
rect 35 -366 39 -357
rect 51 -366 55 -357
rect 18 -370 28 -366
rect 35 -370 44 -366
rect 51 -370 58 -366
rect 76 -366 80 -357
rect 111 -366 115 -357
rect 63 -370 67 -366
rect 76 -370 102 -366
rect 111 -370 125 -366
rect 18 -373 21 -370
rect 35 -373 39 -370
rect 51 -373 55 -370
rect -91 -381 -75 -380
rect -112 -385 -110 -381
rect -103 -384 -75 -381
rect -56 -381 -47 -378
rect -68 -382 -47 -381
rect -40 -382 -24 -378
rect -68 -384 -52 -382
rect -103 -391 -99 -384
rect -68 -391 -64 -384
rect -40 -391 -36 -382
rect -147 -417 -143 -411
rect -111 -417 -107 -411
rect -76 -417 -72 -411
rect -48 -417 -44 -411
rect -143 -421 -137 -417
rect -133 -421 -127 -417
rect -123 -421 -111 -417
rect -107 -421 -103 -417
rect -99 -421 -76 -417
rect -72 -421 -68 -417
rect -64 -421 -48 -417
rect -44 -421 -40 -417
rect -147 -427 -143 -421
rect -111 -427 -107 -421
rect -76 -427 -72 -421
rect -48 -427 -44 -421
rect -27 -436 -24 -382
rect -1 -376 21 -373
rect 60 -377 79 -373
rect -13 -387 -9 -383
rect 27 -387 31 -383
rect 43 -387 47 -383
rect -9 -391 -5 -387
rect -1 -391 27 -387
rect 31 -391 35 -387
rect 39 -391 43 -387
rect 47 -391 51 -387
rect -9 -401 -3 -397
rect 1 -401 7 -397
rect 11 -401 15 -397
rect 19 -401 25 -397
rect 29 -401 33 -397
rect -13 -407 -9 -401
rect 7 -407 11 -401
rect 15 -407 19 -401
rect -3 -436 1 -427
rect 23 -436 27 -427
rect 60 -411 63 -377
rect 86 -380 90 -370
rect 98 -377 114 -373
rect 121 -380 125 -370
rect 125 -400 128 -397
rect 66 -404 70 -400
rect 101 -404 105 -400
rect 70 -408 76 -404
rect 80 -408 86 -404
rect 90 -408 101 -404
rect 105 -408 111 -404
rect 115 -408 121 -404
rect 144 -411 147 -356
rect 159 -363 162 -356
rect 175 -363 178 -349
rect 60 -414 147 -411
rect 181 -349 191 -345
rect 198 -349 207 -345
rect 214 -349 256 -345
rect 263 -349 279 -345
rect 150 -409 154 -403
rect 166 -409 170 -403
rect 181 -409 184 -349
rect 198 -358 202 -349
rect 214 -358 218 -349
rect 254 -358 268 -354
rect 275 -366 279 -349
rect 291 -346 295 -342
rect 326 -346 330 -342
rect 190 -384 194 -378
rect 206 -384 210 -378
rect 194 -388 206 -384
rect 150 -413 184 -409
rect 279 -372 304 -369
rect 311 -375 315 -366
rect 323 -372 339 -369
rect 346 -373 350 -366
rect 354 -352 358 -342
rect 358 -356 362 -352
rect 366 -356 370 -352
rect 374 -356 378 -352
rect 354 -360 358 -356
rect 370 -360 374 -356
rect 362 -373 366 -370
rect 311 -376 327 -375
rect 290 -380 292 -376
rect 299 -379 327 -376
rect 346 -376 355 -373
rect 334 -377 355 -376
rect 362 -377 371 -373
rect 334 -379 350 -377
rect 299 -386 303 -379
rect 334 -386 338 -379
rect 362 -386 366 -377
rect 378 -386 382 -370
rect 255 -412 259 -406
rect 291 -412 295 -406
rect 326 -412 330 -406
rect 354 -412 358 -406
rect 370 -412 374 -406
rect -27 -439 -12 -436
rect -3 -440 16 -436
rect 23 -439 41 -436
rect -36 -447 -21 -444
rect -16 -447 0 -444
rect -112 -457 -110 -453
rect -103 -454 -99 -447
rect -68 -454 -64 -447
rect -103 -457 -75 -454
rect -91 -458 -75 -457
rect -68 -456 -52 -454
rect -68 -457 -47 -456
rect -123 -464 -98 -461
rect -91 -467 -87 -458
rect -56 -460 -47 -457
rect -79 -464 -63 -461
rect -56 -467 -52 -460
rect -40 -463 -36 -447
rect 7 -450 11 -440
rect 23 -443 27 -439
rect -148 -479 -134 -475
rect -127 -484 -123 -467
rect -153 -488 -146 -484
rect -139 -488 -123 -484
rect 15 -457 19 -453
rect 19 -461 25 -457
rect 11 -470 30 -466
rect -48 -477 -44 -473
rect -13 -474 -9 -470
rect -44 -481 -40 -477
rect -9 -478 -3 -474
rect 1 -478 7 -474
rect -139 -491 -135 -488
rect -111 -491 -107 -487
rect -76 -491 -72 -487
rect -48 -491 -44 -481
rect -130 -495 -111 -491
rect -107 -495 -101 -491
rect -97 -495 -91 -491
rect -87 -495 -76 -491
rect -72 -495 -66 -491
rect -62 -495 -56 -491
rect -52 -495 -44 -491
rect -13 -495 21 -491
rect 38 -494 41 -439
rect -147 -505 -143 -501
rect -130 -505 -126 -495
rect -143 -509 -139 -505
rect -135 -509 -126 -505
rect -147 -513 -143 -509
rect -130 -519 -126 -509
rect -13 -501 -9 -495
rect 3 -501 7 -495
rect -130 -523 -111 -519
rect -107 -523 -101 -519
rect -97 -523 -91 -519
rect -87 -523 -76 -519
rect -72 -523 -66 -519
rect -62 -523 -56 -519
rect -52 -523 -44 -519
rect -139 -526 -135 -523
rect -153 -530 -146 -526
rect -139 -530 -123 -526
rect -148 -539 -134 -535
rect -127 -547 -123 -530
rect -111 -527 -107 -523
rect -76 -527 -72 -523
rect -123 -553 -98 -550
rect -91 -556 -87 -547
rect -79 -553 -63 -550
rect -56 -554 -52 -547
rect -48 -533 -44 -523
rect -44 -537 -40 -533
rect -48 -541 -44 -537
rect -4 -548 -1 -541
rect -40 -554 -36 -551
rect -27 -551 4 -548
rect -27 -554 -24 -551
rect -91 -557 -75 -556
rect -112 -561 -110 -557
rect -103 -560 -75 -557
rect -56 -557 -47 -554
rect -68 -558 -47 -557
rect -40 -558 -24 -554
rect -68 -560 -52 -558
rect -103 -567 -99 -560
rect -68 -567 -64 -560
rect -40 -567 -36 -558
rect -147 -593 -143 -587
rect -111 -593 -107 -587
rect -76 -593 -72 -587
rect -48 -593 -44 -587
rect -143 -597 -137 -593
rect -133 -597 -127 -593
rect -123 -597 -111 -593
rect -107 -597 -103 -593
rect -99 -597 -76 -593
rect -72 -597 -68 -593
rect -64 -597 -48 -593
rect -44 -597 -40 -593
rect -147 -603 -143 -597
rect -111 -603 -107 -597
rect -76 -603 -72 -597
rect -48 -603 -44 -597
rect -112 -633 -110 -629
rect -103 -630 -99 -623
rect -68 -630 -64 -623
rect -103 -633 -75 -630
rect -91 -634 -75 -633
rect -68 -632 -52 -630
rect -40 -632 -36 -623
rect -27 -625 -24 -558
rect 12 -555 15 -541
rect -16 -559 -12 -555
rect -8 -559 15 -555
rect 18 -555 21 -495
rect 31 -520 43 -516
rect 27 -526 31 -520
rect 43 -526 47 -520
rect 51 -526 54 -452
rect 60 -512 63 -414
rect 259 -416 265 -412
rect 269 -416 275 -412
rect 279 -416 291 -412
rect 295 -416 299 -412
rect 303 -416 326 -412
rect 330 -416 334 -412
rect 338 -416 354 -412
rect 358 -416 362 -412
rect 366 -416 370 -412
rect 374 -416 378 -412
rect 173 -423 177 -419
rect 181 -423 209 -419
rect 213 -423 217 -419
rect 221 -423 225 -419
rect 229 -423 233 -419
rect 255 -422 259 -416
rect 291 -422 295 -416
rect 326 -422 330 -416
rect 354 -422 358 -416
rect 370 -422 374 -416
rect 169 -427 173 -423
rect 209 -427 213 -423
rect 225 -427 229 -423
rect 181 -437 203 -434
rect 200 -440 203 -437
rect 217 -440 221 -437
rect 233 -440 237 -437
rect 134 -444 170 -441
rect 174 -444 197 -440
rect 163 -448 186 -447
rect 155 -451 186 -448
rect 178 -458 181 -451
rect 194 -458 197 -444
rect 79 -478 86 -474
rect 90 -478 97 -474
rect 101 -478 107 -474
rect 111 -478 129 -474
rect 133 -478 140 -474
rect 144 -478 151 -474
rect 155 -478 161 -474
rect 75 -484 79 -478
rect 97 -484 101 -478
rect 129 -484 133 -478
rect 151 -484 155 -478
rect 85 -513 89 -504
rect 107 -513 111 -504
rect 139 -513 143 -504
rect 161 -513 165 -504
rect 200 -444 210 -440
rect 217 -444 226 -440
rect 233 -444 246 -440
rect 169 -504 173 -498
rect 185 -504 189 -498
rect 200 -504 203 -444
rect 217 -453 221 -444
rect 233 -453 237 -444
rect 209 -479 213 -473
rect 225 -479 229 -473
rect 213 -483 225 -479
rect 243 -479 246 -444
rect 290 -452 292 -448
rect 299 -449 303 -442
rect 334 -449 338 -442
rect 299 -452 327 -449
rect 311 -453 327 -452
rect 334 -451 350 -449
rect 362 -451 366 -442
rect 334 -452 355 -451
rect 279 -459 304 -456
rect 311 -462 315 -453
rect 346 -455 355 -452
rect 362 -455 371 -451
rect 323 -459 339 -456
rect 346 -462 350 -455
rect 362 -458 366 -455
rect 378 -458 382 -442
rect 254 -474 268 -470
rect 275 -479 279 -462
rect 243 -483 256 -479
rect 263 -483 279 -479
rect 354 -472 358 -468
rect 370 -472 374 -468
rect 358 -476 362 -472
rect 366 -476 370 -472
rect 374 -476 378 -472
rect 263 -486 267 -483
rect 291 -486 295 -482
rect 326 -486 330 -482
rect 354 -486 358 -476
rect 272 -490 291 -486
rect 295 -490 301 -486
rect 305 -490 311 -486
rect 315 -490 326 -486
rect 330 -490 336 -486
rect 340 -490 346 -486
rect 350 -490 358 -486
rect 255 -500 259 -496
rect 272 -500 276 -490
rect 259 -504 263 -500
rect 267 -504 276 -500
rect 169 -508 203 -504
rect 65 -517 76 -513
rect 85 -517 130 -513
rect 139 -517 165 -513
rect 87 -524 88 -520
rect 35 -555 39 -546
rect 51 -555 55 -546
rect 63 -531 100 -528
rect 63 -555 66 -531
rect 107 -534 111 -517
rect 18 -559 28 -555
rect 35 -559 44 -555
rect 51 -558 66 -555
rect 18 -562 21 -559
rect 35 -562 39 -559
rect 51 -562 55 -558
rect -1 -565 21 -562
rect -13 -576 -9 -572
rect 27 -576 31 -572
rect 43 -576 47 -572
rect 61 -559 66 -558
rect 51 -576 54 -572
rect -9 -580 -5 -576
rect -1 -580 27 -576
rect 31 -580 35 -576
rect 39 -580 43 -576
rect -9 -590 -3 -586
rect 1 -590 7 -586
rect 11 -590 15 -586
rect 19 -590 23 -586
rect -13 -596 -9 -590
rect 7 -596 11 -590
rect 15 -596 19 -590
rect -3 -625 1 -616
rect 23 -625 27 -616
rect 61 -624 64 -559
rect 115 -524 142 -520
rect 75 -568 79 -564
rect 79 -572 85 -568
rect 89 -572 97 -568
rect 101 -572 107 -568
rect 79 -582 85 -578
rect 89 -582 95 -578
rect 75 -588 79 -582
rect 95 -588 99 -582
rect 72 -617 75 -611
rect 85 -617 89 -608
rect 115 -617 118 -524
rect 72 -621 76 -617
rect 85 -621 118 -617
rect 122 -531 154 -527
rect -27 -628 -12 -625
rect -3 -629 16 -625
rect -68 -633 -47 -632
rect -123 -640 -98 -637
rect -91 -643 -87 -634
rect -56 -636 -47 -633
rect -40 -636 -21 -632
rect -16 -636 0 -633
rect -79 -640 -63 -637
rect -56 -643 -52 -636
rect -40 -639 -36 -636
rect 7 -639 11 -629
rect 61 -628 88 -624
rect 23 -632 27 -630
rect 95 -631 99 -621
rect -148 -655 -134 -651
rect -127 -660 -123 -643
rect -153 -664 -146 -660
rect -139 -664 -123 -660
rect -48 -653 -44 -649
rect -44 -657 -40 -653
rect -139 -667 -135 -664
rect -111 -667 -107 -663
rect -76 -667 -72 -663
rect -48 -667 -44 -657
rect 15 -646 19 -642
rect 19 -650 25 -646
rect 75 -655 79 -651
rect 11 -659 34 -656
rect 79 -659 85 -655
rect 89 -659 95 -655
rect -13 -663 -9 -659
rect 31 -662 34 -659
rect 122 -662 125 -531
rect 161 -534 165 -517
rect 257 -542 261 -538
rect 265 -542 274 -538
rect 253 -546 257 -542
rect 270 -552 274 -542
rect 270 -556 289 -552
rect 293 -556 299 -552
rect 303 -556 309 -552
rect 313 -556 324 -552
rect 328 -556 334 -552
rect 338 -556 344 -552
rect 348 -556 356 -552
rect 261 -559 265 -556
rect 165 -564 171 -561
rect 129 -568 133 -564
rect 133 -572 139 -568
rect 143 -572 151 -568
rect 155 -572 161 -568
rect 168 -575 171 -564
rect -9 -667 -3 -663
rect 1 -667 7 -663
rect 31 -665 125 -662
rect 145 -578 171 -575
rect 233 -563 254 -559
rect 261 -563 277 -559
rect 145 -667 148 -578
rect 155 -650 159 -646
rect 163 -650 191 -646
rect 195 -650 199 -646
rect 203 -650 207 -646
rect 211 -650 215 -646
rect 151 -654 155 -650
rect 191 -654 195 -650
rect 207 -654 211 -650
rect 163 -664 185 -661
rect 182 -667 185 -664
rect 199 -667 203 -664
rect 215 -667 219 -664
rect 233 -667 236 -563
rect 252 -572 266 -568
rect 273 -580 277 -563
rect 289 -560 293 -556
rect 324 -560 328 -556
rect -130 -671 -111 -667
rect -107 -671 -101 -667
rect -97 -671 -91 -667
rect -87 -671 -76 -667
rect -72 -671 -66 -667
rect -62 -671 -56 -667
rect -52 -671 -44 -667
rect 74 -671 138 -668
rect 145 -671 152 -667
rect 156 -671 179 -667
rect -147 -681 -143 -677
rect -130 -681 -126 -671
rect -143 -685 -139 -681
rect -135 -685 -126 -681
rect 74 -713 77 -671
rect 135 -674 138 -671
rect 85 -678 92 -674
rect 96 -678 103 -674
rect 107 -678 114 -674
rect 118 -678 125 -674
rect 135 -678 168 -674
rect 81 -684 85 -678
rect 103 -684 107 -678
rect 125 -684 129 -678
rect 160 -685 163 -678
rect 176 -685 179 -671
rect 91 -707 95 -704
rect 115 -707 119 -704
rect 91 -710 119 -707
rect 52 -716 82 -713
rect -13 -731 21 -727
rect -13 -737 -9 -731
rect 3 -737 7 -731
rect -143 -746 -139 -742
rect -135 -746 -126 -742
rect -147 -750 -143 -746
rect -130 -756 -126 -746
rect -130 -760 -111 -756
rect -107 -760 -101 -756
rect -97 -760 -91 -756
rect -87 -760 -76 -756
rect -72 -760 -66 -756
rect -62 -760 -56 -756
rect -52 -760 -44 -756
rect -139 -763 -135 -760
rect -153 -767 -146 -763
rect -139 -767 -123 -763
rect -148 -776 -134 -772
rect -127 -784 -123 -767
rect -111 -764 -107 -760
rect -76 -764 -72 -760
rect -123 -790 -98 -787
rect -91 -793 -87 -784
rect -79 -790 -63 -787
rect -56 -791 -52 -784
rect -48 -770 -44 -760
rect -44 -774 -40 -770
rect -48 -778 -44 -774
rect -4 -784 -1 -777
rect -40 -791 -36 -788
rect -27 -787 4 -784
rect -27 -791 -24 -787
rect -91 -794 -75 -793
rect -112 -798 -110 -794
rect -103 -797 -75 -794
rect -56 -794 -47 -791
rect -68 -795 -47 -794
rect -40 -795 -24 -791
rect 12 -791 15 -777
rect -16 -795 -12 -791
rect -8 -795 15 -791
rect 18 -791 21 -731
rect 31 -756 43 -752
rect 27 -762 31 -756
rect 43 -762 47 -756
rect 52 -762 55 -716
rect 115 -720 119 -710
rect 79 -724 94 -720
rect 115 -724 129 -720
rect 63 -731 106 -728
rect 72 -738 118 -735
rect 35 -791 39 -782
rect 51 -791 55 -782
rect 18 -795 28 -791
rect 35 -795 44 -791
rect 51 -795 61 -791
rect -68 -797 -52 -795
rect -103 -804 -99 -797
rect -68 -804 -64 -797
rect -40 -804 -36 -795
rect -147 -830 -143 -824
rect -111 -830 -107 -824
rect -76 -830 -72 -824
rect -48 -830 -44 -824
rect -143 -834 -137 -830
rect -133 -834 -127 -830
rect -123 -834 -111 -830
rect -107 -834 -103 -830
rect -99 -834 -76 -830
rect -72 -834 -68 -830
rect -64 -834 -48 -830
rect -44 -834 -40 -830
rect -147 -840 -143 -834
rect -111 -840 -107 -834
rect -76 -840 -72 -834
rect -48 -840 -44 -834
rect -112 -870 -110 -866
rect -103 -867 -99 -860
rect -68 -867 -64 -860
rect -103 -870 -75 -867
rect -91 -871 -75 -870
rect -68 -869 -52 -867
rect -40 -868 -36 -860
rect -27 -861 -24 -795
rect 18 -798 21 -795
rect 35 -798 39 -795
rect 51 -798 55 -795
rect -1 -801 21 -798
rect -13 -812 -9 -808
rect 27 -812 31 -808
rect 43 -812 47 -808
rect -9 -816 -5 -812
rect -1 -816 27 -812
rect 31 -816 35 -812
rect 39 -816 43 -812
rect 47 -816 51 -812
rect -9 -826 -3 -822
rect 1 -826 7 -822
rect 11 -826 15 -822
rect 19 -826 25 -822
rect 29 -826 33 -822
rect -13 -832 -9 -826
rect 7 -832 11 -826
rect 15 -832 19 -826
rect 58 -848 61 -795
rect 75 -833 78 -738
rect 125 -741 129 -724
rect 182 -671 192 -667
rect 199 -671 208 -667
rect 215 -671 236 -667
rect 277 -586 302 -583
rect 309 -589 313 -580
rect 321 -586 337 -583
rect 344 -587 348 -580
rect 352 -566 356 -556
rect 356 -570 360 -566
rect 364 -570 368 -566
rect 372 -570 376 -566
rect 352 -574 356 -570
rect 368 -574 372 -570
rect 360 -587 364 -584
rect 309 -590 325 -589
rect 288 -594 290 -590
rect 297 -593 325 -590
rect 344 -590 353 -587
rect 332 -591 353 -590
rect 360 -591 369 -587
rect 332 -593 348 -591
rect 297 -600 301 -593
rect 332 -600 336 -593
rect 360 -600 364 -591
rect 376 -600 380 -584
rect 253 -626 257 -620
rect 289 -626 293 -620
rect 324 -626 328 -620
rect 352 -626 356 -620
rect 368 -626 372 -620
rect 257 -630 263 -626
rect 267 -630 273 -626
rect 277 -630 289 -626
rect 293 -630 297 -626
rect 301 -630 324 -626
rect 328 -630 332 -626
rect 336 -630 352 -626
rect 356 -630 360 -626
rect 364 -630 368 -626
rect 372 -630 376 -626
rect 253 -636 257 -630
rect 289 -636 293 -630
rect 324 -636 328 -630
rect 352 -636 356 -630
rect 368 -636 372 -630
rect 151 -731 155 -725
rect 167 -731 171 -725
rect 182 -731 185 -671
rect 199 -680 203 -671
rect 215 -680 219 -671
rect 288 -666 290 -662
rect 297 -663 301 -656
rect 332 -663 336 -656
rect 297 -666 325 -663
rect 309 -667 325 -666
rect 332 -665 348 -663
rect 360 -665 364 -656
rect 332 -666 353 -665
rect 277 -673 302 -670
rect 309 -676 313 -667
rect 344 -669 353 -666
rect 360 -669 369 -665
rect 321 -673 337 -670
rect 344 -676 348 -669
rect 360 -672 364 -669
rect 376 -672 380 -656
rect 252 -688 266 -684
rect 273 -693 277 -676
rect 247 -697 254 -693
rect 261 -697 277 -693
rect 352 -686 356 -682
rect 368 -686 372 -682
rect 356 -690 360 -686
rect 364 -690 368 -686
rect 372 -690 376 -686
rect 191 -706 195 -700
rect 207 -706 211 -700
rect 195 -710 207 -706
rect 247 -721 250 -697
rect 261 -700 265 -697
rect 289 -700 293 -696
rect 324 -700 328 -696
rect 352 -700 356 -690
rect 270 -704 289 -700
rect 293 -704 299 -700
rect 303 -704 309 -700
rect 313 -704 324 -700
rect 328 -704 334 -700
rect 338 -704 344 -700
rect 348 -704 356 -700
rect 253 -714 257 -710
rect 270 -714 274 -704
rect 257 -718 261 -714
rect 265 -718 274 -714
rect 247 -724 298 -721
rect 151 -735 185 -731
rect 227 -736 231 -732
rect 235 -736 263 -732
rect 267 -736 271 -732
rect 275 -736 279 -732
rect 283 -736 287 -732
rect 155 -742 162 -738
rect 166 -742 173 -738
rect 177 -742 184 -738
rect 188 -742 195 -738
rect 151 -748 155 -742
rect 173 -748 177 -742
rect 195 -748 199 -742
rect 223 -740 227 -736
rect 263 -740 267 -736
rect 279 -740 283 -736
rect 235 -750 257 -747
rect 254 -753 257 -750
rect 271 -753 275 -750
rect 287 -753 291 -750
rect 295 -753 298 -724
rect 203 -757 224 -753
rect 228 -757 251 -753
rect 161 -771 165 -768
rect 185 -771 189 -768
rect 161 -774 189 -771
rect 129 -781 152 -777
rect 81 -785 85 -781
rect 185 -784 189 -774
rect 203 -784 206 -757
rect 212 -764 240 -760
rect 85 -789 91 -785
rect 95 -789 103 -785
rect 107 -789 115 -785
rect 119 -789 125 -785
rect 132 -788 164 -784
rect 185 -788 199 -784
rect 91 -799 98 -795
rect 102 -799 109 -795
rect 113 -799 119 -795
rect 87 -805 91 -799
rect 109 -805 113 -799
rect 75 -838 76 -833
rect 97 -834 101 -825
rect 119 -834 123 -825
rect 81 -838 88 -834
rect 97 -838 123 -834
rect 119 -841 123 -838
rect 132 -841 135 -788
rect 72 -845 100 -841
rect 119 -845 135 -841
rect 138 -795 176 -791
rect 195 -792 199 -788
rect 212 -792 215 -764
rect 232 -771 235 -764
rect 248 -771 251 -757
rect 195 -795 215 -792
rect 58 -852 112 -848
rect -3 -861 1 -852
rect 23 -861 27 -852
rect -27 -864 -12 -861
rect -3 -865 16 -861
rect -68 -870 -47 -869
rect -123 -877 -98 -874
rect -91 -880 -87 -871
rect -56 -873 -47 -870
rect -40 -872 -21 -868
rect -16 -872 0 -869
rect -79 -877 -63 -874
rect -56 -880 -52 -873
rect -40 -876 -36 -872
rect 7 -875 11 -865
rect 23 -866 28 -861
rect 23 -868 27 -866
rect -148 -892 -134 -888
rect -127 -897 -123 -880
rect -153 -901 -146 -897
rect -139 -901 -123 -897
rect -48 -890 -44 -886
rect -44 -894 -40 -890
rect -139 -904 -135 -901
rect -111 -904 -107 -900
rect -76 -904 -72 -900
rect -48 -904 -44 -894
rect 15 -882 19 -878
rect 19 -886 25 -882
rect 11 -895 57 -892
rect -13 -899 -9 -895
rect -9 -903 -3 -899
rect 1 -903 7 -899
rect -130 -908 -111 -904
rect -107 -908 -101 -904
rect -97 -908 -91 -904
rect -87 -908 -76 -904
rect -72 -908 -66 -904
rect -62 -908 -56 -904
rect -52 -908 -44 -904
rect -147 -918 -143 -914
rect -130 -918 -126 -908
rect -143 -922 -139 -918
rect -135 -922 -126 -918
rect -147 -926 -143 -922
rect -130 -932 -126 -922
rect -130 -936 -111 -932
rect -107 -936 -101 -932
rect -97 -936 -91 -932
rect -87 -936 -76 -932
rect -72 -936 -66 -932
rect -62 -936 -56 -932
rect -52 -936 -44 -932
rect -139 -939 -135 -936
rect -153 -943 -146 -939
rect -139 -943 -123 -939
rect -148 -952 -134 -948
rect -127 -960 -123 -943
rect -111 -940 -107 -936
rect -76 -940 -72 -936
rect -123 -966 -98 -963
rect -91 -969 -87 -960
rect -79 -966 -63 -963
rect -56 -967 -52 -960
rect -48 -946 -44 -936
rect -44 -950 -40 -946
rect -48 -954 -44 -950
rect -91 -970 -75 -969
rect -112 -974 -110 -970
rect -103 -973 -75 -970
rect -56 -970 -47 -967
rect -68 -971 -47 -970
rect -68 -973 -52 -971
rect -103 -980 -99 -973
rect -68 -980 -64 -973
rect -40 -980 -36 -964
rect 54 -983 57 -895
rect 76 -936 79 -852
rect 119 -855 123 -845
rect 87 -889 91 -885
rect 91 -893 98 -889
rect 102 -893 108 -889
rect 112 -893 119 -889
rect 91 -903 97 -899
rect 101 -903 107 -899
rect 87 -909 91 -903
rect 107 -909 111 -903
rect 75 -938 79 -936
rect 97 -938 101 -929
rect 138 -938 141 -795
rect 75 -941 88 -938
rect 97 -942 141 -938
rect 144 -802 188 -798
rect 78 -949 100 -945
rect 107 -952 111 -942
rect 144 -945 148 -802
rect 195 -805 199 -795
rect 254 -757 264 -753
rect 271 -757 280 -753
rect 287 -757 298 -753
rect 223 -817 227 -811
rect 239 -817 243 -811
rect 254 -817 257 -757
rect 271 -766 275 -757
rect 287 -766 291 -757
rect 263 -792 267 -786
rect 279 -792 283 -786
rect 267 -796 279 -792
rect 223 -821 257 -817
rect 151 -849 155 -845
rect 155 -853 161 -849
rect 165 -853 173 -849
rect 177 -853 185 -849
rect 189 -853 195 -849
rect 114 -948 148 -945
rect 87 -976 91 -972
rect 91 -980 97 -976
rect 101 -980 107 -976
rect 114 -983 117 -948
rect 54 -986 117 -983
rect -36 -1000 48 -996
rect 79 -998 86 -994
rect 90 -998 97 -994
rect 101 -998 108 -994
rect 112 -998 121 -994
rect 125 -998 131 -994
rect -147 -1006 -143 -1000
rect -111 -1006 -107 -1000
rect -76 -1006 -72 -1000
rect -48 -1006 -44 -1000
rect 75 -1004 79 -998
rect 97 -1004 101 -998
rect 121 -1004 125 -998
rect -143 -1010 -137 -1006
rect -133 -1010 -127 -1006
rect -123 -1010 -111 -1006
rect -107 -1010 -103 -1006
rect -99 -1010 -76 -1006
rect -72 -1010 -68 -1006
rect -64 -1010 -48 -1006
rect -44 -1010 -40 -1006
rect 85 -1027 89 -1024
rect 109 -1027 113 -1024
rect 131 -1027 135 -1024
rect 85 -1030 135 -1027
rect 71 -1037 76 -1033
rect 68 -1042 88 -1040
rect 63 -1044 88 -1042
rect 60 -1051 100 -1047
rect 72 -1058 112 -1054
rect 121 -1062 124 -1051
rect 58 -1065 124 -1062
rect -13 -1112 21 -1108
rect -13 -1118 -9 -1112
rect 3 -1118 7 -1112
rect -143 -1127 -139 -1123
rect -135 -1127 -126 -1123
rect -147 -1131 -143 -1127
rect -130 -1137 -126 -1127
rect -130 -1141 -111 -1137
rect -107 -1141 -101 -1137
rect -97 -1141 -91 -1137
rect -87 -1141 -76 -1137
rect -72 -1141 -66 -1137
rect -62 -1141 -56 -1137
rect -52 -1141 -44 -1137
rect -139 -1144 -135 -1141
rect -153 -1148 -146 -1144
rect -139 -1148 -123 -1144
rect -148 -1157 -134 -1153
rect -127 -1165 -123 -1148
rect -111 -1145 -107 -1141
rect -76 -1145 -72 -1141
rect -123 -1171 -98 -1168
rect -91 -1174 -87 -1165
rect -79 -1171 -63 -1168
rect -56 -1172 -52 -1165
rect -48 -1151 -44 -1141
rect -44 -1155 -40 -1151
rect -48 -1159 -44 -1155
rect -4 -1165 -1 -1158
rect -40 -1172 -36 -1169
rect -27 -1168 4 -1165
rect -27 -1172 -24 -1168
rect -91 -1175 -75 -1174
rect -112 -1179 -110 -1175
rect -103 -1178 -75 -1175
rect -56 -1175 -47 -1172
rect -68 -1176 -47 -1175
rect -40 -1176 -24 -1172
rect 12 -1172 15 -1158
rect -16 -1176 -12 -1172
rect -8 -1176 15 -1172
rect 18 -1172 21 -1112
rect 31 -1137 43 -1133
rect 27 -1143 31 -1137
rect 43 -1143 47 -1137
rect 35 -1172 39 -1163
rect 51 -1172 55 -1163
rect 58 -1172 61 -1065
rect 131 -1068 135 -1030
rect 135 -1118 141 -1115
rect 75 -1122 79 -1118
rect 79 -1126 85 -1122
rect 89 -1126 97 -1122
rect 101 -1126 109 -1122
rect 113 -1126 121 -1122
rect 125 -1126 131 -1122
rect 87 -1138 94 -1134
rect 98 -1138 105 -1134
rect 109 -1138 116 -1134
rect 120 -1138 127 -1134
rect 83 -1144 87 -1138
rect 105 -1144 109 -1138
rect 127 -1144 131 -1138
rect 93 -1167 97 -1164
rect 117 -1167 121 -1164
rect 93 -1170 121 -1167
rect 18 -1176 28 -1172
rect 35 -1176 44 -1172
rect 51 -1176 61 -1172
rect -68 -1178 -52 -1176
rect -103 -1185 -99 -1178
rect -68 -1185 -64 -1178
rect -40 -1185 -36 -1176
rect -147 -1211 -143 -1205
rect -111 -1211 -107 -1205
rect -76 -1211 -72 -1205
rect -48 -1211 -44 -1205
rect -143 -1215 -137 -1211
rect -133 -1215 -127 -1211
rect -123 -1215 -111 -1211
rect -107 -1215 -103 -1211
rect -99 -1215 -76 -1211
rect -72 -1215 -68 -1211
rect -64 -1215 -48 -1211
rect -44 -1215 -40 -1211
rect -147 -1221 -143 -1215
rect -111 -1221 -107 -1215
rect -76 -1221 -72 -1215
rect -48 -1221 -44 -1215
rect -112 -1251 -110 -1247
rect -103 -1248 -99 -1241
rect -68 -1248 -64 -1241
rect -103 -1251 -75 -1248
rect -91 -1252 -75 -1251
rect -68 -1250 -52 -1248
rect -40 -1249 -36 -1241
rect -27 -1242 -24 -1176
rect 18 -1179 21 -1176
rect 35 -1179 39 -1176
rect 51 -1179 55 -1176
rect -1 -1182 21 -1179
rect 58 -1187 61 -1176
rect 78 -1176 84 -1173
rect 117 -1180 121 -1170
rect 138 -1173 141 -1118
rect 226 -1124 232 -1120
rect 236 -1124 242 -1120
rect 246 -1124 258 -1120
rect 262 -1124 266 -1120
rect 270 -1124 293 -1120
rect 297 -1124 301 -1120
rect 305 -1124 321 -1120
rect 325 -1124 329 -1120
rect 333 -1124 337 -1120
rect 341 -1124 345 -1120
rect 222 -1130 226 -1124
rect 258 -1130 262 -1124
rect 293 -1130 297 -1124
rect 321 -1130 325 -1124
rect 337 -1130 341 -1124
rect 158 -1138 165 -1134
rect 169 -1138 176 -1134
rect 180 -1138 187 -1134
rect 191 -1138 200 -1134
rect 204 -1138 210 -1134
rect 154 -1144 158 -1138
rect 176 -1144 180 -1138
rect 200 -1144 204 -1138
rect 164 -1167 168 -1164
rect 188 -1167 192 -1164
rect 210 -1167 214 -1164
rect 164 -1170 214 -1167
rect 257 -1160 259 -1156
rect 266 -1157 270 -1150
rect 301 -1157 305 -1150
rect 266 -1160 294 -1157
rect 278 -1161 294 -1160
rect 301 -1159 317 -1157
rect 329 -1159 333 -1150
rect 301 -1160 322 -1159
rect 246 -1167 271 -1164
rect 278 -1170 282 -1161
rect 313 -1163 322 -1160
rect 329 -1163 338 -1159
rect 290 -1167 306 -1164
rect 313 -1170 317 -1163
rect 329 -1166 333 -1163
rect 345 -1166 349 -1150
rect 138 -1177 155 -1173
rect 69 -1184 96 -1181
rect 117 -1184 167 -1180
rect -13 -1193 -9 -1189
rect 27 -1193 31 -1189
rect 43 -1193 47 -1189
rect 58 -1190 108 -1187
rect -9 -1197 -5 -1193
rect -1 -1197 27 -1193
rect 31 -1197 35 -1193
rect 39 -1197 43 -1193
rect 47 -1197 51 -1193
rect -9 -1207 -3 -1203
rect 1 -1207 7 -1203
rect 11 -1207 15 -1203
rect 19 -1207 25 -1203
rect 29 -1207 33 -1203
rect -13 -1213 -9 -1207
rect 7 -1213 11 -1207
rect 15 -1213 19 -1207
rect -3 -1242 1 -1233
rect -27 -1245 -12 -1242
rect -3 -1246 16 -1242
rect -68 -1251 -47 -1250
rect -123 -1258 -98 -1255
rect -91 -1261 -87 -1252
rect -56 -1254 -47 -1251
rect -40 -1253 -21 -1249
rect -16 -1253 0 -1250
rect -79 -1258 -63 -1255
rect -56 -1261 -52 -1254
rect -40 -1257 -36 -1253
rect 7 -1256 11 -1246
rect 23 -1249 27 -1233
rect -148 -1273 -134 -1269
rect -127 -1278 -123 -1261
rect -153 -1282 -146 -1278
rect -139 -1282 -123 -1278
rect -48 -1271 -44 -1267
rect -44 -1275 -40 -1271
rect -139 -1285 -135 -1282
rect -111 -1285 -107 -1281
rect -76 -1285 -72 -1281
rect -48 -1285 -44 -1275
rect 15 -1263 19 -1259
rect 19 -1267 25 -1263
rect 32 -1272 35 -1256
rect 11 -1276 35 -1272
rect -13 -1280 -9 -1276
rect -9 -1284 -3 -1280
rect 1 -1284 7 -1280
rect -130 -1289 -111 -1285
rect -107 -1289 -101 -1285
rect -97 -1289 -91 -1285
rect -87 -1289 -76 -1285
rect -72 -1289 -66 -1285
rect -62 -1289 -56 -1285
rect -52 -1289 -44 -1285
rect -147 -1299 -143 -1295
rect -130 -1299 -126 -1289
rect -143 -1303 -139 -1299
rect -135 -1303 -126 -1299
rect 58 -1310 61 -1190
rect 98 -1198 120 -1195
rect 127 -1201 131 -1184
rect 210 -1187 214 -1170
rect 225 -1182 235 -1178
rect 242 -1187 246 -1170
rect 134 -1191 179 -1187
rect 210 -1191 223 -1187
rect 230 -1191 246 -1187
rect 321 -1180 325 -1176
rect 337 -1180 341 -1176
rect 325 -1184 329 -1180
rect 333 -1184 337 -1180
rect 341 -1184 345 -1180
rect 83 -1245 87 -1241
rect 87 -1249 93 -1245
rect 97 -1249 105 -1245
rect 109 -1249 117 -1245
rect 121 -1249 127 -1245
rect 97 -1261 104 -1257
rect 108 -1261 115 -1257
rect 119 -1261 125 -1257
rect 93 -1267 97 -1261
rect 115 -1267 119 -1261
rect 134 -1267 137 -1191
rect 129 -1270 137 -1267
rect 140 -1198 191 -1194
rect 84 -1296 86 -1295
rect 103 -1296 107 -1287
rect 125 -1296 129 -1287
rect 84 -1298 94 -1296
rect 82 -1300 94 -1298
rect 103 -1300 129 -1296
rect 78 -1307 106 -1303
rect 58 -1314 118 -1310
rect 87 -1401 90 -1314
rect 125 -1317 129 -1300
rect 93 -1351 97 -1347
rect 97 -1355 104 -1351
rect 108 -1355 114 -1351
rect 118 -1355 125 -1351
rect 107 -1366 113 -1362
rect 117 -1366 123 -1362
rect 103 -1372 107 -1366
rect 123 -1372 127 -1366
rect 113 -1401 117 -1392
rect 140 -1401 143 -1198
rect 147 -1205 203 -1201
rect 147 -1249 150 -1205
rect 210 -1208 214 -1191
rect 230 -1194 234 -1191
rect 258 -1194 262 -1190
rect 293 -1194 297 -1190
rect 321 -1194 325 -1184
rect 239 -1198 258 -1194
rect 262 -1198 268 -1194
rect 272 -1198 293 -1194
rect 297 -1198 303 -1194
rect 307 -1198 313 -1194
rect 317 -1198 325 -1194
rect 222 -1208 226 -1204
rect 239 -1208 243 -1198
rect 226 -1212 230 -1208
rect 234 -1212 243 -1208
rect 154 -1262 158 -1258
rect 158 -1266 164 -1262
rect 168 -1266 176 -1262
rect 180 -1266 188 -1262
rect 192 -1266 200 -1262
rect 204 -1266 210 -1262
rect 87 -1405 104 -1401
rect 113 -1405 143 -1401
rect 86 -1412 116 -1408
rect 123 -1415 127 -1405
rect 103 -1439 107 -1435
rect 107 -1443 113 -1439
rect 117 -1443 123 -1439
<< m2contact >>
rect 85 -21 90 -16
rect 118 -29 123 -24
rect 53 -43 58 -38
rect -153 -363 -148 -358
rect -84 -377 -79 -372
rect -21 -370 -16 -365
rect -117 -385 -112 -380
rect 93 -378 98 -373
rect 249 -358 254 -353
rect 318 -372 323 -367
rect 285 -380 290 -375
rect -21 -447 -16 -442
rect -117 -458 -112 -453
rect -84 -466 -79 -461
rect -153 -480 -148 -475
rect 30 -470 35 -465
rect 50 -452 55 -447
rect -153 -539 -148 -534
rect -84 -553 -79 -548
rect -117 -561 -112 -556
rect -117 -634 -112 -629
rect -21 -559 -16 -554
rect 150 -452 155 -447
rect 60 -517 65 -512
rect 285 -453 290 -448
rect 318 -461 323 -456
rect 249 -475 254 -470
rect 50 -581 55 -576
rect -21 -636 -16 -631
rect -84 -642 -79 -637
rect 23 -630 28 -625
rect -153 -656 -148 -651
rect 247 -572 252 -567
rect -153 -776 -148 -771
rect -84 -790 -79 -785
rect -117 -798 -112 -793
rect -21 -795 -16 -790
rect 74 -724 79 -719
rect 67 -740 72 -735
rect -117 -871 -112 -866
rect 316 -586 321 -581
rect 283 -594 288 -589
rect 283 -667 288 -662
rect 316 -675 321 -670
rect 247 -689 252 -684
rect -21 -872 -16 -867
rect -84 -879 -79 -874
rect -153 -893 -148 -888
rect -153 -952 -148 -947
rect -84 -966 -79 -961
rect -117 -974 -112 -969
rect 73 -950 78 -945
rect 48 -1000 53 -995
rect 67 -1059 72 -1054
rect -153 -1157 -148 -1152
rect -84 -1171 -79 -1166
rect -117 -1179 -112 -1174
rect -21 -1176 -16 -1171
rect -117 -1252 -112 -1247
rect 252 -1161 257 -1156
rect 285 -1169 290 -1164
rect -21 -1253 -16 -1248
rect -84 -1260 -79 -1255
rect -153 -1274 -148 -1269
rect 220 -1183 225 -1178
rect 79 -1298 84 -1293
<< metal2 >>
rect 85 -26 89 -21
rect 85 -29 118 -26
rect 85 -43 89 -29
rect 53 -46 89 -43
rect -19 -299 27 -296
rect -19 -337 -16 -299
rect 24 -320 27 -299
rect 24 -324 252 -320
rect -82 -340 -16 -337
rect -153 -366 -113 -363
rect -153 -475 -150 -366
rect -117 -372 -113 -366
rect -82 -372 -79 -340
rect 249 -353 252 -324
rect 249 -361 289 -358
rect -117 -375 -84 -372
rect -117 -380 -113 -375
rect -19 -442 -16 -370
rect 94 -409 97 -378
rect 31 -412 97 -409
rect -117 -463 -113 -458
rect -117 -466 -84 -463
rect 31 -465 34 -412
rect 55 -451 150 -448
rect -117 -480 -113 -466
rect 249 -467 252 -361
rect 285 -367 289 -361
rect 285 -370 318 -367
rect 285 -375 289 -370
rect 285 -458 289 -453
rect 285 -461 318 -458
rect 285 -467 289 -461
rect 249 -470 289 -467
rect -153 -483 -113 -480
rect -153 -531 -150 -483
rect 37 -508 42 -503
rect -153 -534 -113 -531
rect -153 -651 -150 -539
rect -117 -548 -113 -534
rect -117 -551 -84 -548
rect -117 -556 -113 -551
rect -19 -631 -16 -559
rect 28 -629 46 -626
rect -117 -639 -113 -634
rect -117 -642 -84 -639
rect -117 -656 -113 -642
rect -153 -659 -113 -656
rect -153 -768 -150 -659
rect 43 -744 46 -629
rect 51 -737 54 -581
rect 60 -720 63 -517
rect 249 -532 252 -475
rect 247 -535 252 -532
rect 247 -567 250 -535
rect 67 -574 72 -569
rect 247 -575 287 -572
rect 247 -681 250 -575
rect 283 -581 287 -575
rect 283 -584 316 -581
rect 283 -589 287 -584
rect 283 -672 287 -667
rect 283 -675 316 -672
rect 283 -681 287 -675
rect 247 -684 287 -681
rect 60 -723 74 -720
rect 51 -740 67 -737
rect 43 -747 63 -744
rect -153 -771 -113 -768
rect -153 -888 -150 -776
rect -117 -785 -113 -771
rect -117 -788 -84 -785
rect -117 -793 -113 -788
rect -19 -867 -16 -795
rect -117 -876 -113 -871
rect -117 -879 -84 -876
rect -117 -893 -113 -879
rect -153 -896 -113 -893
rect -153 -944 -150 -896
rect -153 -947 -113 -944
rect 60 -945 63 -747
rect 76 -826 79 -724
rect 317 -822 320 -675
rect 286 -825 320 -822
rect 76 -829 88 -826
rect 85 -851 88 -829
rect 82 -854 88 -851
rect 60 -946 73 -945
rect -153 -1149 -150 -952
rect -117 -961 -113 -947
rect 41 -949 73 -946
rect -117 -964 -84 -961
rect -117 -969 -113 -964
rect 41 -1066 44 -949
rect 82 -987 85 -854
rect 48 -990 85 -987
rect 48 -995 51 -990
rect 48 -1055 51 -1000
rect 48 -1058 67 -1055
rect 41 -1069 59 -1066
rect -153 -1152 -113 -1149
rect -153 -1269 -150 -1157
rect -117 -1166 -113 -1152
rect -117 -1169 -84 -1166
rect -117 -1174 -113 -1169
rect -19 -1248 -16 -1176
rect -117 -1257 -113 -1252
rect -117 -1260 -84 -1257
rect -117 -1274 -113 -1260
rect -153 -1277 -113 -1274
rect 56 -1294 59 -1069
rect 252 -1166 256 -1161
rect 286 -1164 289 -825
rect 252 -1169 285 -1166
rect 252 -1183 256 -1169
rect 220 -1186 256 -1183
rect 56 -1298 79 -1294
<< m3contact >>
rect 23 -866 28 -861
<< m123contact >>
rect 132 -349 137 -344
rect 58 -370 63 -365
rect 128 -402 133 -397
rect 129 -444 134 -439
rect 37 -499 42 -494
rect 82 -525 87 -520
rect 67 -614 72 -609
rect 58 -733 63 -728
rect 202 -789 207 -784
rect 76 -838 81 -833
rect 67 -845 72 -840
rect 70 -941 75 -936
rect 70 -1033 75 -1028
rect 63 -1042 68 -1037
rect 55 -1051 60 -1046
rect 120 -1051 125 -1046
rect 31 -1256 36 -1251
rect 73 -1177 78 -1172
rect 64 -1184 69 -1179
rect 93 -1198 98 -1193
rect 146 -1254 151 -1249
rect 73 -1307 78 -1302
rect 81 -1413 86 -1408
<< metal3 >>
rect 128 -349 132 -345
rect 128 -362 131 -349
rect 59 -365 131 -362
rect 38 -503 41 -499
rect 58 -521 61 -370
rect 129 -439 132 -402
rect 58 -525 82 -521
rect 58 -728 61 -525
rect 68 -609 71 -574
rect 28 -865 38 -862
rect 35 -1072 38 -865
rect 59 -920 62 -733
rect 68 -840 71 -614
rect 68 -855 71 -845
rect 56 -923 62 -920
rect 56 -1046 59 -923
rect 78 -928 81 -838
rect 203 -856 206 -789
rect 63 -931 81 -928
rect 151 -859 206 -856
rect 63 -1037 66 -931
rect 70 -1028 73 -941
rect 151 -951 154 -859
rect 140 -954 154 -951
rect 35 -1075 60 -1072
rect 36 -1255 40 -1252
rect 57 -1317 60 -1075
rect 64 -1179 67 -1042
rect 72 -1046 75 -1033
rect 71 -1049 75 -1046
rect 71 -1128 74 -1049
rect 140 -1047 143 -954
rect 125 -1050 143 -1047
rect 71 -1131 76 -1128
rect 73 -1172 76 -1131
rect 73 -1302 76 -1177
rect 85 -1198 93 -1195
rect 85 -1254 146 -1251
rect 57 -1320 84 -1317
rect 81 -1408 84 -1320
<< m345contact >>
rect 37 -508 42 -503
rect 67 -574 72 -569
rect 67 -860 72 -855
rect 80 -1198 85 -1193
rect 40 -1256 45 -1251
rect 80 -1256 85 -1251
<< metal5 >>
rect 42 -507 71 -504
rect 68 -569 71 -507
rect 68 -1195 71 -860
rect 68 -1198 80 -1195
rect 45 -1255 80 -1252
<< labels >>
rlabel metal1 93 -476 93 -476 1 vdd
rlabel metal1 55 -368 55 -368 1 p0
rlabel metal1 123 -368 123 -368 1 c1
rlabel metal1 22 -468 22 -468 1 g0_inv
rlabel metal1 25 -438 25 -438 1 g0
rlabel metal1 118 -329 118 -329 1 vdd
rlabel metal1 83 -329 83 -329 1 vdd
rlabel metal1 83 -406 83 -406 1 gnd
rlabel metal2 -18 -373 -18 -373 1 b0
rlabel metal1 -25 -361 -25 -361 1 a0
rlabel metal1 22 -459 22 -459 1 gnd
rlabel metal1 4 -476 4 -476 1 gnd
rlabel metal1 4 -399 4 -399 1 vdd
rlabel metal1 13 -389 13 -389 1 gnd
rlabel metal1 37 -329 37 -329 1 vdd
rlabel metal1 53 -557 53 -557 1 p1
rlabel metal1 22 -648 22 -648 1 gnd
rlabel metal1 4 -665 4 -665 1 gnd
rlabel metal1 4 -588 4 -588 1 vdd
rlabel metal1 13 -578 13 -578 1 gnd
rlabel metal1 37 -518 37 -518 1 vdd
rlabel metal1 25 -624 25 -624 1 g1
rlabel metal1 93 -570 93 -570 1 gnd
rlabel metal1 147 -570 147 -570 1 gnd
rlabel metal1 92 -580 92 -580 1 vdd
rlabel metal1 92 -657 92 -657 1 gnd
rlabel metal1 13 -658 13 -658 1 g1_inv
rlabel metal1 -14 -51 -14 -51 1 gnd
rlabel metal1 304 -182 304 -182 7 out_NAND5
rlabel metal1 236 -196 236 -196 1 in5_NAND5
rlabel metal1 236 -189 236 -189 1 in4_NAND5
rlabel metal1 236 -182 236 -182 1 in3_NAND5
rlabel metal1 236 -175 236 -175 1 in2_NAND5
rlabel metal1 236 -168 236 -168 1 in1_NAND5
rlabel metal1 258 -257 258 -257 1 gnd
rlabel metal1 257 -129 257 -129 1 vdd
rlabel space 122 -246 190 -120 1 NAND4
rlabel metal1 184 -175 184 -175 7 out_NAND4
rlabel metal1 128 -189 128 -189 1 in4_NAND4
rlabel metal1 128 -182 128 -182 1 in3_NAND4
rlabel metal1 128 -175 128 -175 1 in2_NAND4
rlabel metal1 128 -168 128 -168 1 in1_NAND4
rlabel metal1 150 -240 150 -240 1 gnd
rlabel metal1 149 -129 149 -129 1 vdd
rlabel space 47 -230 104 -117 1 NAND3
rlabel metal1 98 -175 98 -175 7 out_NAND3
rlabel metal1 76 -223 76 -223 1 gnd
rlabel metal1 76 -129 76 -129 1 vdd
rlabel metal1 54 -182 54 -182 1 in3_NAND3
rlabel metal1 54 -175 54 -175 1 in2_NAND3
rlabel metal1 54 -168 54 -168 1 in1_NAND3
rlabel metal1 15 -168 15 -168 1 out_NAND2
rlabel metal1 4 -206 4 -206 1 gnd
rlabel metal1 -17 -175 -17 -175 1 in2_NAND2
rlabel metal1 -17 -168 -17 -168 1 in1_NAND2
rlabel metal1 4 -129 4 -129 1 vdd
rlabel space -23 -216 28 -119 1 NAND2
rlabel metal1 262 -6 262 -6 1 vdd
rlabel metal1 284 -45 284 -45 1 out_xor
rlabel metal1 208 -45 208 -45 1 in1_xor
rlabel metal1 208 -38 208 -38 1 in2_xor
rlabel space 202 -79 293 29 1 xor
rlabel metal1 238 -66 238 -66 1 gnd
rlabel metal1 -14 9 -14 9 1 vdd
rlabel metal1 -4 -30 -4 -30 1 out_inv
rlabel metal1 -24 -30 -24 -30 1 in_inv
rlabel metal1 170 -21 170 -21 1 out_ff
rlabel metal1 51 -40 51 -40 1 clk
rlabel metal1 51 -49 51 -49 1 in_ff
rlabel space 46 -75 177 26 1 flipflop
rlabel space -33 -60 3 19 1 inverter
rlabel metal1 195 -421 195 -421 5 gnd
rlabel metal1 200 -386 200 -386 5 vdd
rlabel metal1 176 -326 176 -326 5 gnd
rlabel metal1 171 -1136 171 -1136 1 vdd
rlabel metal1 172 -1264 172 -1264 1 gnd
rlabel metal1 25 -1244 25 -1244 1 g3
rlabel metal1 13 -1274 13 -1274 1 g3_inv
rlabel metal1 25 -860 25 -860 1 g2
rlabel metal1 120 -1441 120 -1441 1 gnd
rlabel metal1 120 -1364 120 -1364 1 vdd
rlabel metal1 53 -1174 53 -1174 1 p3
rlabel metal1 111 -1353 111 -1353 1 gnd
rlabel metal1 111 -1259 111 -1259 1 vdd
rlabel metal1 101 -1247 101 -1247 1 gnd
rlabel metal1 100 -1136 100 -1136 1 vdd
rlabel metal1 53 -793 53 -793 1 p2
rlabel metal1 93 -1124 93 -1124 1 gnd
rlabel metal1 92 -996 92 -996 1 vdd
rlabel metal1 169 -851 169 -851 1 gnd
rlabel metal1 168 -740 168 -740 1 vdd
rlabel metal1 13 -894 13 -894 1 g2_inv
rlabel metal1 37 -754 37 -754 1 vdd
rlabel metal1 13 -814 13 -814 1 gnd
rlabel metal1 4 -824 4 -824 1 vdd
rlabel metal1 4 -901 4 -901 1 gnd
rlabel metal1 22 -884 22 -884 1 gnd
rlabel metal1 98 -676 98 -676 1 vdd
rlabel metal1 99 -787 99 -787 1 gnd
rlabel metal1 105 -797 105 -797 1 vdd
rlabel metal1 105 -891 105 -891 1 gnd
rlabel metal1 104 -978 104 -978 1 gnd
rlabel metal1 104 -901 104 -901 1 vdd
rlabel metal1 37 -1135 37 -1135 1 vdd
rlabel metal1 13 -1195 13 -1195 1 gnd
rlabel metal1 4 -1205 4 -1205 1 vdd
rlabel metal1 4 -1282 4 -1282 1 gnd
rlabel metal1 22 -1265 22 -1265 1 gnd
rlabel metal1 163 -522 163 -522 1 c2
rlabel metal1 177 -648 177 -648 5 gnd
rlabel metal1 201 -708 201 -708 5 vdd
rlabel metal1 197 -786 197 -786 1 c3
rlabel metal1 -151 -352 -151 -352 3 a0_ff_in
rlabel metal1 -82 -669 -82 -669 1 gnd
rlabel metal1 -128 -507 -128 -507 1 gnd
rlabel metal1 -151 -486 -151 -486 3 b0_ff_in
rlabel metal1 -31 -556 -31 -556 1 a1
rlabel metal1 -151 -528 -151 -528 3 a1_ff_in
rlabel metal1 -151 -662 -151 -662 3 b1_ff_in
rlabel metal1 -28 -634 -28 -634 1 b1
rlabel metal1 112 18 112 18 1 vdd
rlabel metal1 115 -56 115 -56 1 gnd
rlabel metal1 -128 -920 -128 -920 1 gnd
rlabel metal1 -82 -758 -82 -758 1 gnd
rlabel metal1 -28 -870 -28 -870 1 b2
rlabel metal1 -28 -793 -28 -793 1 a2
rlabel metal1 -151 -941 -151 -941 3 c0_ff_in
rlabel metal1 -88 -832 -88 -832 1 vdd
rlabel metal1 -87 -1008 -87 -1008 1 vdd
rlabel metal1 30 -998 30 -998 1 c0
rlabel metal1 -88 -1213 -88 -1213 1 vdd
rlabel metal1 -82 -1139 -82 -1139 1 gnd
rlabel metal1 -128 -1301 -128 -1301 1 gnd
rlabel metal1 -28 -1174 -28 -1174 1 a3
rlabel metal1 -28 -1251 -28 -1251 1 b3
rlabel metal1 -151 -1280 -151 -1280 3 b3_ff_in
rlabel metal1 -151 -1146 -151 -1146 3 a3_ff_in
rlabel metal1 -151 -765 -151 -765 3 a2_ff_in
rlabel metal1 -151 -899 -151 -899 3 b2_ff_in
rlabel metal1 320 -340 320 -340 1 gnd
rlabel metal1 274 -502 274 -502 1 gnd
rlabel metal1 237 -347 237 -347 1 s0
rlabel metal1 364 -375 364 -375 1 s0_ff_out
rlabel metal1 364 -452 364 -452 1 s1_ff_out
rlabel metal1 244 -442 244 -442 1 s1
rlabel metal1 -88 -419 -88 -419 1 vdd
rlabel metal1 -87 -595 -87 -595 1 vdd
rlabel metal1 318 -554 318 -554 1 gnd
rlabel metal1 272 -716 272 -716 1 gnd
rlabel metal1 311 -628 311 -628 1 vdd
rlabel metal1 314 -414 314 -414 1 vdd
rlabel metal1 228 -669 228 -669 1 s2
rlabel metal1 -84 -345 -84 -345 1 gnd
rlabel metal1 279 -1122 279 -1122 1 vdd
rlabel metal1 282 -1196 282 -1196 1 gnd
rlabel metal1 212 -1189 212 -1189 1 c4
rlabel metal2 -151 -364 -151 -364 3 clk
rlabel metal1 362 -589 362 -589 1 s2_ff_out
rlabel metal1 362 -666 362 -666 1 s3_ff_out
rlabel metal1 337 -1161 337 -1161 1 c4_ff_out
rlabel metal1 380 -375 380 -375 1 s0_ff_out_inv
rlabel metal1 380 -453 380 -453 1 s1_ff_out_inv
rlabel metal1 378 -589 378 -589 1 s2_ff_out_inv
rlabel metal1 378 -667 378 -667 1 s3_ff_out_inv
rlabel metal1 347 -1161 347 -1161 1 c4_ff_out_inv
rlabel metal1 249 -734 249 -734 5 gnd
rlabel metal1 273 -794 273 -794 5 vdd
rlabel metal1 289 -755 289 -755 1 s3
<< end >>
