magic
tech scmos
timestamp 1731862927
<< nwell >>
rect -26 -25 -2 14
rect 49 -16 172 23
rect 206 -1 246 24
rect 49 -36 85 -16
rect 206 -35 286 -1
rect 246 -40 286 -35
rect -19 -163 17 -124
rect 52 -163 100 -124
rect 126 -163 186 -124
rect 234 -163 306 -124
rect -19 -331 21 -306
rect -19 -365 61 -331
rect 21 -370 61 -365
rect -19 -440 33 -401
rect -19 -513 21 -488
rect -19 -547 61 -513
rect 21 -552 61 -547
rect -19 -622 33 -583
rect -19 -697 21 -672
rect -19 -731 61 -697
rect 21 -736 61 -731
rect -19 -806 33 -767
rect -19 -879 21 -854
rect -19 -913 61 -879
rect 21 -918 61 -913
rect -19 -988 33 -949
<< ntransistor >>
rect -15 -45 -13 -35
rect 96 -50 98 -30
rect 108 -50 110 -30
rect 131 -50 133 -30
rect 143 -50 145 -30
rect 159 -36 161 -26
rect 60 -64 62 -54
rect 217 -60 219 -50
rect 257 -60 259 -50
rect 273 -60 275 -50
rect -8 -200 -6 -180
rect 4 -200 6 -180
rect 63 -217 65 -187
rect 75 -217 77 -187
rect 87 -217 89 -187
rect 137 -234 139 -194
rect 149 -234 151 -194
rect 161 -234 163 -194
rect 173 -234 175 -194
rect 245 -251 247 -201
rect 257 -251 259 -201
rect 269 -251 271 -201
rect 281 -251 283 -201
rect 293 -251 295 -201
rect -8 -390 -6 -380
rect 32 -390 34 -380
rect 48 -390 50 -380
rect -8 -477 -6 -457
rect 4 -477 6 -457
rect 20 -460 22 -450
rect -8 -572 -6 -562
rect 32 -572 34 -562
rect 48 -572 50 -562
rect -8 -659 -6 -639
rect 4 -659 6 -639
rect 20 -642 22 -632
rect -8 -756 -6 -746
rect 32 -756 34 -746
rect 48 -756 50 -746
rect -8 -843 -6 -823
rect 4 -843 6 -823
rect 20 -826 22 -816
rect -8 -938 -6 -928
rect 32 -938 34 -928
rect 48 -938 50 -928
rect -8 -1025 -6 -1005
rect 4 -1025 6 -1005
rect 20 -1008 22 -998
<< ptransistor >>
rect -15 -19 -13 1
rect 60 -30 62 10
rect 72 -30 74 10
rect 96 -10 98 10
rect 131 -10 133 10
rect 159 -10 161 10
rect 217 -29 219 11
rect 233 -29 235 11
rect 257 -34 259 -14
rect 273 -34 275 -14
rect -8 -157 -6 -137
rect 4 -157 6 -137
rect 63 -157 65 -137
rect 75 -157 77 -137
rect 87 -157 89 -137
rect 137 -157 139 -137
rect 149 -157 151 -137
rect 161 -157 163 -137
rect 173 -157 175 -137
rect 245 -157 247 -137
rect 257 -157 259 -137
rect 269 -157 271 -137
rect 281 -157 283 -137
rect 293 -157 295 -137
rect -8 -359 -6 -319
rect 8 -359 10 -319
rect 32 -364 34 -344
rect 48 -364 50 -344
rect -8 -434 -6 -414
rect 4 -434 6 -414
rect 20 -434 22 -414
rect -8 -541 -6 -501
rect 8 -541 10 -501
rect 32 -546 34 -526
rect 48 -546 50 -526
rect -8 -616 -6 -596
rect 4 -616 6 -596
rect 20 -616 22 -596
rect -8 -725 -6 -685
rect 8 -725 10 -685
rect 32 -730 34 -710
rect 48 -730 50 -710
rect -8 -800 -6 -780
rect 4 -800 6 -780
rect 20 -800 22 -780
rect -8 -907 -6 -867
rect 8 -907 10 -867
rect 32 -912 34 -892
rect 48 -912 50 -892
rect -8 -982 -6 -962
rect 4 -982 6 -962
rect 20 -982 22 -962
<< ndiffusion >>
rect -16 -45 -15 -35
rect -13 -45 -12 -35
rect 95 -50 96 -30
rect 98 -50 108 -30
rect 110 -50 111 -30
rect 130 -50 131 -30
rect 133 -50 143 -30
rect 145 -50 146 -30
rect 158 -36 159 -26
rect 161 -36 162 -26
rect 59 -64 60 -54
rect 62 -64 63 -54
rect 216 -60 217 -50
rect 219 -60 220 -50
rect 256 -60 257 -50
rect 259 -60 260 -50
rect 272 -60 273 -50
rect 275 -60 276 -50
rect -9 -200 -8 -180
rect -6 -200 4 -180
rect 6 -200 7 -180
rect 62 -217 63 -187
rect 65 -217 75 -187
rect 77 -217 87 -187
rect 89 -217 90 -187
rect 136 -234 137 -194
rect 139 -234 149 -194
rect 151 -234 161 -194
rect 163 -234 173 -194
rect 175 -234 176 -194
rect 244 -251 245 -201
rect 247 -251 257 -201
rect 259 -251 269 -201
rect 271 -251 281 -201
rect 283 -251 293 -201
rect 295 -251 296 -201
rect -9 -390 -8 -380
rect -6 -390 -5 -380
rect 31 -390 32 -380
rect 34 -390 35 -380
rect 47 -390 48 -380
rect 50 -390 51 -380
rect -9 -477 -8 -457
rect -6 -477 4 -457
rect 6 -477 7 -457
rect 19 -460 20 -450
rect 22 -460 23 -450
rect -9 -572 -8 -562
rect -6 -572 -5 -562
rect 31 -572 32 -562
rect 34 -572 35 -562
rect 47 -572 48 -562
rect 50 -572 51 -562
rect -9 -659 -8 -639
rect -6 -659 4 -639
rect 6 -659 7 -639
rect 19 -642 20 -632
rect 22 -642 23 -632
rect -9 -756 -8 -746
rect -6 -756 -5 -746
rect 31 -756 32 -746
rect 34 -756 35 -746
rect 47 -756 48 -746
rect 50 -756 51 -746
rect -9 -843 -8 -823
rect -6 -843 4 -823
rect 6 -843 7 -823
rect 19 -826 20 -816
rect 22 -826 23 -816
rect -9 -938 -8 -928
rect -6 -938 -5 -928
rect 31 -938 32 -928
rect 34 -938 35 -928
rect 47 -938 48 -928
rect 50 -938 51 -928
rect -9 -1025 -8 -1005
rect -6 -1025 4 -1005
rect 6 -1025 7 -1005
rect 19 -1008 20 -998
rect 22 -1008 23 -998
<< pdiffusion >>
rect -16 -19 -15 1
rect -13 -19 -12 1
rect 59 -30 60 10
rect 62 -30 72 10
rect 74 -30 75 10
rect 95 -10 96 10
rect 98 -10 99 10
rect 130 -10 131 10
rect 133 -10 134 10
rect 158 -10 159 10
rect 161 -10 162 10
rect 216 -29 217 11
rect 219 -29 220 11
rect 232 -29 233 11
rect 235 -29 236 11
rect 256 -34 257 -14
rect 259 -34 260 -14
rect 272 -34 273 -14
rect 275 -34 276 -14
rect -9 -157 -8 -137
rect -6 -157 -5 -137
rect 3 -157 4 -137
rect 6 -157 7 -137
rect 62 -157 63 -137
rect 65 -157 66 -137
rect 74 -157 75 -137
rect 77 -157 78 -137
rect 86 -157 87 -137
rect 89 -157 90 -137
rect 136 -157 137 -137
rect 139 -157 140 -137
rect 148 -157 149 -137
rect 151 -157 152 -137
rect 160 -157 161 -137
rect 163 -157 164 -137
rect 172 -157 173 -137
rect 175 -157 176 -137
rect 244 -157 245 -137
rect 247 -157 248 -137
rect 256 -157 257 -137
rect 259 -157 260 -137
rect 268 -157 269 -137
rect 271 -157 272 -137
rect 280 -157 281 -137
rect 283 -157 284 -137
rect 292 -157 293 -137
rect 295 -157 296 -137
rect -9 -359 -8 -319
rect -6 -359 -5 -319
rect 7 -359 8 -319
rect 10 -359 11 -319
rect 31 -364 32 -344
rect 34 -364 35 -344
rect 47 -364 48 -344
rect 50 -364 51 -344
rect -9 -434 -8 -414
rect -6 -434 -5 -414
rect 3 -434 4 -414
rect 6 -434 7 -414
rect 19 -434 20 -414
rect 22 -434 23 -414
rect -9 -541 -8 -501
rect -6 -541 -5 -501
rect 7 -541 8 -501
rect 10 -541 11 -501
rect 31 -546 32 -526
rect 34 -546 35 -526
rect 47 -546 48 -526
rect 50 -546 51 -526
rect -9 -616 -8 -596
rect -6 -616 -5 -596
rect 3 -616 4 -596
rect 6 -616 7 -596
rect 19 -616 20 -596
rect 22 -616 23 -596
rect -9 -725 -8 -685
rect -6 -725 -5 -685
rect 7 -725 8 -685
rect 10 -725 11 -685
rect 31 -730 32 -710
rect 34 -730 35 -710
rect 47 -730 48 -710
rect 50 -730 51 -710
rect -9 -800 -8 -780
rect -6 -800 -5 -780
rect 3 -800 4 -780
rect 6 -800 7 -780
rect 19 -800 20 -780
rect 22 -800 23 -780
rect -9 -907 -8 -867
rect -6 -907 -5 -867
rect 7 -907 8 -867
rect 10 -907 11 -867
rect 31 -912 32 -892
rect 34 -912 35 -892
rect 47 -912 48 -892
rect 50 -912 51 -892
rect -9 -982 -8 -962
rect -6 -982 -5 -962
rect 3 -982 4 -962
rect 6 -982 7 -962
rect 19 -982 20 -962
rect 22 -982 23 -962
<< ndcontact >>
rect -20 -45 -16 -35
rect -12 -45 -8 -35
rect 91 -50 95 -30
rect 111 -50 115 -30
rect 126 -50 130 -30
rect 146 -50 150 -30
rect 154 -36 158 -26
rect 162 -36 166 -26
rect 55 -64 59 -54
rect 63 -64 67 -54
rect 212 -60 216 -50
rect 220 -60 224 -50
rect 252 -60 256 -50
rect 260 -60 264 -50
rect 268 -60 272 -50
rect 276 -60 280 -50
rect -13 -200 -9 -180
rect 7 -200 11 -180
rect 58 -217 62 -187
rect 90 -217 94 -187
rect 132 -234 136 -194
rect 176 -234 180 -194
rect 240 -251 244 -201
rect 296 -251 300 -201
rect -13 -390 -9 -380
rect -5 -390 -1 -380
rect 27 -390 31 -380
rect 35 -390 39 -380
rect 43 -390 47 -380
rect 51 -390 55 -380
rect -13 -477 -9 -457
rect 7 -477 11 -457
rect 15 -460 19 -450
rect 23 -460 27 -450
rect -13 -572 -9 -562
rect -5 -572 -1 -562
rect 27 -572 31 -562
rect 35 -572 39 -562
rect 43 -572 47 -562
rect 51 -572 55 -562
rect -13 -659 -9 -639
rect 7 -659 11 -639
rect 15 -642 19 -632
rect 23 -642 27 -632
rect -13 -756 -9 -746
rect -5 -756 -1 -746
rect 27 -756 31 -746
rect 35 -756 39 -746
rect 43 -756 47 -746
rect 51 -756 55 -746
rect -13 -843 -9 -823
rect 7 -843 11 -823
rect 15 -826 19 -816
rect 23 -826 27 -816
rect -13 -938 -9 -928
rect -5 -938 -1 -928
rect 27 -938 31 -928
rect 35 -938 39 -928
rect 43 -938 47 -928
rect 51 -938 55 -928
rect -13 -1025 -9 -1005
rect 7 -1025 11 -1005
rect 15 -1008 19 -998
rect 23 -1008 27 -998
<< pdcontact >>
rect -20 -19 -16 1
rect -12 -19 -8 1
rect 55 -30 59 10
rect 75 -30 79 10
rect 91 -10 95 10
rect 99 -10 103 10
rect 126 -10 130 10
rect 134 -10 138 10
rect 154 -10 158 10
rect 162 -10 166 10
rect 212 -29 216 11
rect 220 -29 224 11
rect 228 -29 232 11
rect 236 -29 240 11
rect 252 -34 256 -14
rect 260 -34 264 -14
rect 268 -34 272 -14
rect 276 -34 280 -14
rect -13 -157 -9 -137
rect -5 -157 3 -137
rect 7 -157 11 -137
rect 58 -157 62 -137
rect 66 -157 74 -137
rect 78 -157 86 -137
rect 90 -157 94 -137
rect 132 -157 136 -137
rect 140 -157 148 -137
rect 152 -157 160 -137
rect 164 -157 172 -137
rect 176 -157 180 -137
rect 240 -157 244 -137
rect 248 -157 256 -137
rect 260 -157 268 -137
rect 272 -157 280 -137
rect 284 -157 292 -137
rect 296 -157 300 -137
rect -13 -359 -9 -319
rect -5 -359 -1 -319
rect 3 -359 7 -319
rect 11 -359 15 -319
rect 27 -364 31 -344
rect 35 -364 39 -344
rect 43 -364 47 -344
rect 51 -364 55 -344
rect -13 -434 -9 -414
rect -5 -434 3 -414
rect 7 -434 11 -414
rect 15 -434 19 -414
rect 23 -434 27 -414
rect -13 -541 -9 -501
rect -5 -541 -1 -501
rect 3 -541 7 -501
rect 11 -541 15 -501
rect 27 -546 31 -526
rect 35 -546 39 -526
rect 43 -546 47 -526
rect 51 -546 55 -526
rect -13 -616 -9 -596
rect -5 -616 3 -596
rect 7 -616 11 -596
rect 15 -616 19 -596
rect 23 -616 27 -596
rect -13 -725 -9 -685
rect -5 -725 -1 -685
rect 3 -725 7 -685
rect 11 -725 15 -685
rect 27 -730 31 -710
rect 35 -730 39 -710
rect 43 -730 47 -710
rect 51 -730 55 -710
rect -13 -800 -9 -780
rect -5 -800 3 -780
rect 7 -800 11 -780
rect 15 -800 19 -780
rect 23 -800 27 -780
rect -13 -907 -9 -867
rect -5 -907 -1 -867
rect 3 -907 7 -867
rect 11 -907 15 -867
rect 27 -912 31 -892
rect 35 -912 39 -892
rect 43 -912 47 -892
rect 51 -912 55 -892
rect -13 -982 -9 -962
rect -5 -982 3 -962
rect 7 -982 11 -962
rect 15 -982 19 -962
rect 23 -982 27 -962
<< psubstratepcontact >>
rect -20 -53 -16 -49
rect -12 -53 -8 -49
rect 154 -44 158 -40
rect 164 -44 168 -40
rect 72 -58 76 -54
rect 87 -58 91 -54
rect 103 -58 107 -54
rect 122 -58 126 -54
rect 138 -58 142 -54
rect 154 -58 158 -54
rect 212 -68 216 -64
rect 220 -68 224 -64
rect 252 -68 256 -64
rect 260 -68 264 -64
rect 268 -68 272 -64
rect 276 -68 280 -64
rect 51 -72 55 -68
rect 62 -72 66 -68
rect 72 -72 76 -68
rect -13 -208 -9 -204
rect -3 -208 1 -204
rect 7 -208 11 -204
rect 58 -225 62 -221
rect 69 -225 73 -221
rect 79 -225 83 -221
rect 90 -225 94 -221
rect 132 -242 136 -238
rect 142 -242 146 -238
rect 154 -242 158 -238
rect 166 -242 170 -238
rect 176 -242 180 -238
rect 240 -259 244 -255
rect 250 -259 254 -255
rect 262 -259 266 -255
rect 274 -259 278 -255
rect 286 -259 290 -255
rect 296 -259 300 -255
rect -13 -398 -9 -394
rect -5 -398 -1 -394
rect 27 -398 31 -394
rect 35 -398 39 -394
rect 43 -398 47 -394
rect 51 -398 55 -394
rect 15 -468 19 -464
rect 25 -468 29 -464
rect -13 -485 -9 -481
rect -3 -485 1 -481
rect 7 -485 11 -481
rect -13 -580 -9 -576
rect -5 -580 -1 -576
rect 27 -580 31 -576
rect 35 -580 39 -576
rect 43 -580 47 -576
rect 51 -580 55 -576
rect 15 -650 19 -646
rect 25 -650 29 -646
rect -13 -667 -9 -663
rect -3 -667 1 -663
rect 7 -667 11 -663
rect -13 -764 -9 -760
rect -5 -764 -1 -760
rect 27 -764 31 -760
rect 35 -764 39 -760
rect 43 -764 47 -760
rect 51 -764 55 -760
rect 15 -834 19 -830
rect 25 -834 29 -830
rect -13 -851 -9 -847
rect -3 -851 1 -847
rect 7 -851 11 -847
rect -13 -946 -9 -942
rect -5 -946 -1 -942
rect 27 -946 31 -942
rect 35 -946 39 -942
rect 43 -946 47 -942
rect 51 -946 55 -942
rect 15 -1016 19 -1012
rect 25 -1016 29 -1012
rect -13 -1033 -9 -1029
rect -3 -1033 1 -1029
rect 7 -1033 11 -1029
<< nsubstratencontact >>
rect 53 16 57 20
rect 65 16 69 20
rect 76 16 80 20
rect 87 16 91 20
rect 101 16 105 20
rect 112 16 116 20
rect 122 16 126 20
rect 136 16 140 20
rect 152 16 156 20
rect 164 16 168 20
rect -20 7 -16 11
rect -12 7 -8 11
rect 252 -8 256 -4
rect 268 -8 272 -4
rect -13 -131 -9 -127
rect -3 -131 1 -127
rect 7 -131 11 -127
rect 58 -131 62 -127
rect 69 -131 73 -127
rect 80 -131 84 -127
rect 90 -131 94 -127
rect 132 -131 136 -127
rect 143 -131 147 -127
rect 154 -131 158 -127
rect 165 -131 169 -127
rect 176 -131 180 -127
rect 240 -131 244 -127
rect 251 -131 255 -127
rect 262 -131 266 -127
rect 273 -131 277 -127
rect 286 -131 290 -127
rect 296 -131 300 -127
rect 27 -338 31 -334
rect 43 -338 47 -334
rect -13 -408 -9 -404
rect -3 -408 1 -404
rect 7 -408 11 -404
rect 15 -408 19 -404
rect 25 -408 29 -404
rect 27 -520 31 -516
rect 43 -520 47 -516
rect -13 -590 -9 -586
rect -3 -590 1 -586
rect 7 -590 11 -586
rect 15 -590 19 -586
rect 25 -590 29 -586
rect 27 -704 31 -700
rect 43 -704 47 -700
rect -13 -774 -9 -770
rect -3 -774 1 -770
rect 7 -774 11 -770
rect 15 -774 19 -770
rect 25 -774 29 -770
rect 27 -886 31 -882
rect 43 -886 47 -882
rect -13 -956 -9 -952
rect -3 -956 1 -952
rect 7 -956 11 -952
rect 15 -956 19 -952
rect 25 -956 29 -952
<< polysilicon >>
rect 60 10 62 13
rect 72 10 74 13
rect 96 10 98 13
rect 131 10 133 13
rect 159 10 161 13
rect 217 11 219 14
rect 233 11 235 14
rect -15 1 -13 4
rect -15 -35 -13 -19
rect 96 -30 98 -10
rect 108 -30 110 -23
rect 131 -30 133 -10
rect 143 -30 145 -23
rect 159 -26 161 -10
rect -15 -48 -13 -45
rect 60 -54 62 -30
rect 72 -44 74 -30
rect 257 -14 259 -11
rect 273 -14 275 -11
rect 159 -39 161 -36
rect 217 -50 219 -29
rect 233 -40 235 -29
rect 257 -50 259 -34
rect 273 -50 275 -34
rect 96 -53 98 -50
rect 108 -53 110 -50
rect 131 -53 133 -50
rect 143 -53 145 -50
rect 217 -63 219 -60
rect 257 -63 259 -60
rect 273 -63 275 -60
rect 60 -67 62 -64
rect -8 -137 -6 -134
rect 4 -137 6 -134
rect 63 -137 65 -134
rect 75 -137 77 -134
rect 87 -137 89 -134
rect 137 -137 139 -134
rect 149 -137 151 -134
rect 161 -137 163 -134
rect 173 -137 175 -134
rect 245 -137 247 -134
rect 257 -137 259 -134
rect 269 -137 271 -134
rect 281 -137 283 -134
rect 293 -137 295 -134
rect -8 -180 -6 -157
rect 4 -180 6 -157
rect 63 -187 65 -157
rect 75 -187 77 -157
rect 87 -187 89 -157
rect -8 -203 -6 -200
rect 4 -203 6 -200
rect 137 -194 139 -157
rect 149 -194 151 -157
rect 161 -194 163 -157
rect 173 -194 175 -157
rect 63 -220 65 -217
rect 75 -220 77 -217
rect 87 -220 89 -217
rect 245 -201 247 -157
rect 257 -201 259 -157
rect 269 -201 271 -157
rect 281 -201 283 -157
rect 293 -201 295 -157
rect 137 -237 139 -234
rect 149 -237 151 -234
rect 161 -237 163 -234
rect 173 -237 175 -234
rect 245 -254 247 -251
rect 257 -254 259 -251
rect 269 -254 271 -251
rect 281 -254 283 -251
rect 293 -254 295 -251
rect -8 -319 -6 -316
rect 8 -319 10 -316
rect 32 -344 34 -341
rect 48 -344 50 -341
rect -8 -380 -6 -359
rect 8 -370 10 -359
rect 32 -380 34 -364
rect 48 -380 50 -364
rect -8 -393 -6 -390
rect 32 -393 34 -390
rect 48 -393 50 -390
rect -8 -414 -6 -411
rect 4 -414 6 -411
rect 20 -414 22 -411
rect -8 -457 -6 -434
rect 4 -457 6 -434
rect 20 -450 22 -434
rect 20 -463 22 -460
rect -8 -480 -6 -477
rect 4 -480 6 -477
rect -8 -501 -6 -498
rect 8 -501 10 -498
rect 32 -526 34 -523
rect 48 -526 50 -523
rect -8 -562 -6 -541
rect 8 -552 10 -541
rect 32 -562 34 -546
rect 48 -562 50 -546
rect -8 -575 -6 -572
rect 32 -575 34 -572
rect 48 -575 50 -572
rect -8 -596 -6 -593
rect 4 -596 6 -593
rect 20 -596 22 -593
rect -8 -639 -6 -616
rect 4 -639 6 -616
rect 20 -632 22 -616
rect 20 -645 22 -642
rect -8 -662 -6 -659
rect 4 -662 6 -659
rect -8 -685 -6 -682
rect 8 -685 10 -682
rect 32 -710 34 -707
rect 48 -710 50 -707
rect -8 -746 -6 -725
rect 8 -736 10 -725
rect 32 -746 34 -730
rect 48 -746 50 -730
rect -8 -759 -6 -756
rect 32 -759 34 -756
rect 48 -759 50 -756
rect -8 -780 -6 -777
rect 4 -780 6 -777
rect 20 -780 22 -777
rect -8 -823 -6 -800
rect 4 -823 6 -800
rect 20 -816 22 -800
rect 20 -829 22 -826
rect -8 -846 -6 -843
rect 4 -846 6 -843
rect -8 -867 -6 -864
rect 8 -867 10 -864
rect 32 -892 34 -889
rect 48 -892 50 -889
rect -8 -928 -6 -907
rect 8 -918 10 -907
rect 32 -928 34 -912
rect 48 -928 50 -912
rect -8 -941 -6 -938
rect 32 -941 34 -938
rect 48 -941 50 -938
rect -8 -962 -6 -959
rect 4 -962 6 -959
rect 20 -962 22 -959
rect -8 -1005 -6 -982
rect 4 -1005 6 -982
rect 20 -998 22 -982
rect 20 -1011 22 -1008
rect -8 -1028 -6 -1025
rect 4 -1028 6 -1025
<< polycontact >>
rect -19 -32 -15 -28
rect 92 -20 96 -16
rect 127 -21 131 -17
rect 104 -27 108 -23
rect 155 -23 159 -19
rect 139 -27 143 -23
rect 56 -51 60 -47
rect 68 -42 72 -38
rect 213 -47 217 -43
rect 229 -40 233 -36
rect 253 -47 257 -43
rect 269 -47 273 -43
rect -12 -170 -8 -166
rect 0 -177 4 -173
rect 59 -170 63 -166
rect 71 -177 75 -173
rect 83 -184 87 -180
rect 133 -170 137 -166
rect 145 -177 149 -173
rect 157 -184 161 -180
rect 169 -191 173 -187
rect 241 -170 245 -166
rect 253 -177 257 -173
rect 265 -184 269 -180
rect 277 -191 281 -187
rect 289 -198 293 -194
rect -12 -377 -8 -373
rect 4 -370 8 -366
rect 28 -377 32 -373
rect 44 -377 48 -373
rect -12 -447 -8 -443
rect 0 -454 4 -450
rect 16 -447 20 -443
rect -12 -559 -8 -555
rect 4 -552 8 -548
rect 28 -559 32 -555
rect 44 -559 48 -555
rect -12 -629 -8 -625
rect 0 -636 4 -632
rect 16 -629 20 -625
rect -12 -743 -8 -739
rect 4 -736 8 -732
rect 28 -743 32 -739
rect 44 -743 48 -739
rect -12 -813 -8 -809
rect 0 -820 4 -816
rect 16 -813 20 -809
rect -12 -925 -8 -921
rect 4 -918 8 -914
rect 28 -925 32 -921
rect 44 -925 48 -921
rect -12 -995 -8 -991
rect 0 -1002 4 -998
rect 16 -995 20 -991
<< metal1 >>
rect 49 16 53 20
rect 57 16 65 20
rect 69 16 76 20
rect 80 16 87 20
rect 91 16 101 20
rect 105 16 112 20
rect 116 16 122 20
rect 126 16 136 20
rect 140 16 152 20
rect 156 16 164 20
rect 168 16 172 20
rect 212 17 246 21
rect -16 7 -12 11
rect 55 10 59 16
rect 91 10 95 16
rect 126 10 130 16
rect 154 10 158 16
rect 212 11 216 17
rect 228 11 232 17
rect -20 1 -16 7
rect -12 -28 -8 -19
rect -26 -32 -19 -28
rect -12 -32 -2 -28
rect 90 -20 92 -16
rect 99 -17 103 -10
rect 134 -17 138 -10
rect 99 -20 127 -17
rect 111 -21 127 -20
rect 134 -19 150 -17
rect 162 -19 166 -10
rect 134 -20 155 -19
rect 79 -27 104 -24
rect 111 -30 115 -21
rect 146 -23 155 -20
rect 162 -23 172 -19
rect 123 -27 139 -24
rect 146 -30 150 -23
rect 162 -26 166 -23
rect -12 -35 -8 -32
rect 49 -42 53 -38
rect 58 -42 68 -38
rect -20 -49 -16 -45
rect 75 -47 79 -30
rect -16 -53 -12 -49
rect 49 -51 56 -47
rect 63 -51 79 -47
rect 221 -36 224 -29
rect 154 -40 158 -36
rect 206 -40 229 -36
rect 158 -44 164 -40
rect 168 -44 172 -40
rect 237 -43 240 -29
rect 63 -54 67 -51
rect 91 -54 95 -50
rect 126 -54 130 -50
rect 154 -54 158 -44
rect 206 -47 213 -43
rect 217 -47 240 -43
rect 243 -43 246 17
rect 256 -8 268 -4
rect 252 -14 256 -8
rect 268 -14 272 -8
rect 260 -43 264 -34
rect 276 -43 280 -34
rect 243 -47 253 -43
rect 260 -47 269 -43
rect 276 -47 286 -43
rect 243 -50 246 -47
rect 260 -50 264 -47
rect 276 -50 280 -47
rect 76 -58 87 -54
rect 91 -58 103 -54
rect 107 -58 122 -54
rect 126 -58 138 -54
rect 142 -58 154 -54
rect 55 -68 59 -64
rect 72 -68 76 -58
rect 224 -53 246 -50
rect 212 -64 216 -60
rect 252 -64 256 -60
rect 268 -64 272 -60
rect 216 -68 220 -64
rect 224 -68 252 -64
rect 256 -68 260 -64
rect 264 -68 268 -64
rect 272 -68 276 -64
rect 49 -72 51 -68
rect 55 -72 62 -68
rect 66 -72 72 -68
rect -9 -131 -3 -127
rect 1 -131 7 -127
rect -13 -137 -9 -131
rect 7 -137 11 -131
rect 62 -131 69 -127
rect 73 -131 80 -127
rect 84 -131 90 -127
rect 136 -131 143 -127
rect 147 -131 154 -127
rect 158 -131 165 -127
rect 169 -131 176 -127
rect 58 -137 62 -131
rect 80 -137 84 -131
rect 132 -137 136 -131
rect 154 -137 158 -131
rect 176 -137 180 -131
rect 244 -131 251 -127
rect 255 -131 262 -127
rect 266 -131 273 -127
rect 277 -131 286 -127
rect 290 -131 296 -127
rect 240 -137 244 -131
rect 262 -137 266 -131
rect 286 -137 290 -131
rect -3 -166 1 -157
rect 68 -166 72 -157
rect 90 -166 94 -157
rect 142 -160 146 -157
rect 166 -160 170 -157
rect 142 -163 170 -160
rect 250 -160 254 -157
rect 274 -160 278 -157
rect 296 -160 300 -157
rect 250 -163 300 -160
rect -19 -170 -12 -166
rect -3 -170 17 -166
rect 52 -170 59 -166
rect 68 -170 94 -166
rect 126 -170 133 -166
rect -19 -177 0 -173
rect 7 -180 11 -170
rect 90 -173 94 -170
rect 166 -173 170 -163
rect 234 -170 241 -166
rect 52 -177 71 -173
rect 90 -177 100 -173
rect 126 -177 145 -173
rect 166 -177 186 -173
rect 234 -177 253 -173
rect 52 -184 83 -180
rect 90 -187 94 -177
rect 126 -184 157 -180
rect -13 -204 -9 -200
rect -9 -208 -3 -204
rect 1 -208 7 -204
rect 126 -191 169 -187
rect 176 -194 180 -177
rect 296 -180 300 -163
rect 234 -184 265 -180
rect 296 -184 306 -180
rect 234 -191 277 -187
rect 58 -221 62 -217
rect 62 -225 69 -221
rect 73 -225 79 -221
rect 83 -225 90 -221
rect 234 -198 289 -194
rect 296 -201 300 -184
rect 132 -238 136 -234
rect 136 -242 142 -238
rect 146 -242 154 -238
rect 158 -242 166 -238
rect 170 -242 176 -238
rect 240 -255 244 -251
rect 244 -259 250 -255
rect 254 -259 262 -255
rect 266 -259 274 -255
rect 278 -259 286 -255
rect 290 -259 296 -255
rect -13 -313 21 -309
rect -13 -319 -9 -313
rect 3 -319 7 -313
rect -4 -366 -1 -359
rect -27 -369 4 -366
rect -27 -443 -24 -369
rect 12 -373 15 -359
rect -16 -377 -12 -373
rect -8 -377 15 -373
rect 18 -373 21 -313
rect 31 -338 43 -334
rect 27 -344 31 -338
rect 43 -344 47 -338
rect 35 -373 39 -364
rect 51 -373 55 -364
rect 18 -377 28 -373
rect 35 -377 44 -373
rect 51 -377 61 -373
rect 18 -380 21 -377
rect 35 -380 39 -377
rect 51 -380 55 -377
rect -1 -383 21 -380
rect -13 -394 -9 -390
rect 27 -394 31 -390
rect 43 -394 47 -390
rect -9 -398 -5 -394
rect -1 -398 27 -394
rect 31 -398 35 -394
rect 39 -398 43 -394
rect 47 -398 51 -394
rect -9 -408 -3 -404
rect 1 -408 7 -404
rect 11 -408 15 -404
rect 19 -408 25 -404
rect 29 -408 33 -404
rect -13 -414 -9 -408
rect 7 -414 11 -408
rect 15 -414 19 -408
rect -3 -443 1 -434
rect 23 -443 27 -434
rect -27 -446 -12 -443
rect -3 -447 16 -443
rect 23 -447 33 -443
rect -16 -454 0 -451
rect 7 -457 11 -447
rect 23 -450 27 -447
rect 15 -464 19 -460
rect 19 -468 25 -464
rect 11 -477 33 -473
rect -13 -481 -9 -477
rect -9 -485 -3 -481
rect 1 -485 7 -481
rect -13 -495 21 -491
rect -13 -501 -9 -495
rect 3 -501 7 -495
rect -4 -548 -1 -541
rect -27 -551 4 -548
rect -27 -625 -24 -551
rect 12 -555 15 -541
rect -16 -559 -12 -555
rect -8 -559 15 -555
rect 18 -555 21 -495
rect 31 -520 43 -516
rect 27 -526 31 -520
rect 43 -526 47 -520
rect 35 -555 39 -546
rect 51 -555 55 -546
rect 18 -559 28 -555
rect 35 -559 44 -555
rect 51 -559 61 -555
rect 18 -562 21 -559
rect 35 -562 39 -559
rect 51 -562 55 -559
rect -1 -565 21 -562
rect -13 -576 -9 -572
rect 27 -576 31 -572
rect 43 -576 47 -572
rect -9 -580 -5 -576
rect -1 -580 27 -576
rect 31 -580 35 -576
rect 39 -580 43 -576
rect 47 -580 51 -576
rect -9 -590 -3 -586
rect 1 -590 7 -586
rect 11 -590 15 -586
rect 19 -590 25 -586
rect 29 -590 33 -586
rect -13 -596 -9 -590
rect 7 -596 11 -590
rect 15 -596 19 -590
rect -3 -625 1 -616
rect 23 -625 27 -616
rect -27 -628 -12 -625
rect -3 -629 16 -625
rect 23 -629 33 -625
rect -16 -636 0 -633
rect 7 -639 11 -629
rect 23 -632 27 -629
rect 15 -646 19 -642
rect 19 -650 25 -646
rect 11 -659 33 -655
rect -13 -663 -9 -659
rect -9 -667 -3 -663
rect 1 -667 7 -663
rect -13 -679 21 -675
rect -13 -685 -9 -679
rect 3 -685 7 -679
rect -4 -732 -1 -725
rect -27 -735 4 -732
rect -27 -809 -24 -735
rect 12 -739 15 -725
rect -16 -743 -12 -739
rect -8 -743 15 -739
rect 18 -739 21 -679
rect 31 -704 43 -700
rect 27 -710 31 -704
rect 43 -710 47 -704
rect 35 -739 39 -730
rect 51 -739 55 -730
rect 18 -743 28 -739
rect 35 -743 44 -739
rect 51 -743 61 -739
rect 18 -746 21 -743
rect 35 -746 39 -743
rect 51 -746 55 -743
rect -1 -749 21 -746
rect -13 -760 -9 -756
rect 27 -760 31 -756
rect 43 -760 47 -756
rect -9 -764 -5 -760
rect -1 -764 27 -760
rect 31 -764 35 -760
rect 39 -764 43 -760
rect 47 -764 51 -760
rect -9 -774 -3 -770
rect 1 -774 7 -770
rect 11 -774 15 -770
rect 19 -774 25 -770
rect 29 -774 33 -770
rect -13 -780 -9 -774
rect 7 -780 11 -774
rect 15 -780 19 -774
rect -3 -809 1 -800
rect 23 -809 27 -800
rect -27 -812 -12 -809
rect -3 -813 16 -809
rect 23 -813 33 -809
rect -16 -820 0 -817
rect 7 -823 11 -813
rect 23 -816 27 -813
rect 15 -830 19 -826
rect 19 -834 25 -830
rect 11 -843 33 -839
rect -13 -847 -9 -843
rect -9 -851 -3 -847
rect 1 -851 7 -847
rect -13 -861 21 -857
rect -13 -867 -9 -861
rect 3 -867 7 -861
rect -4 -914 -1 -907
rect -27 -917 4 -914
rect -27 -991 -24 -917
rect 12 -921 15 -907
rect -16 -925 -12 -921
rect -8 -925 15 -921
rect 18 -921 21 -861
rect 31 -886 43 -882
rect 27 -892 31 -886
rect 43 -892 47 -886
rect 35 -921 39 -912
rect 51 -921 55 -912
rect 18 -925 28 -921
rect 35 -925 44 -921
rect 51 -925 61 -921
rect 18 -928 21 -925
rect 35 -928 39 -925
rect 51 -928 55 -925
rect -1 -931 21 -928
rect -13 -942 -9 -938
rect 27 -942 31 -938
rect 43 -942 47 -938
rect -9 -946 -5 -942
rect -1 -946 27 -942
rect 31 -946 35 -942
rect 39 -946 43 -942
rect 47 -946 51 -942
rect -9 -956 -3 -952
rect 1 -956 7 -952
rect 11 -956 15 -952
rect 19 -956 25 -952
rect 29 -956 33 -952
rect -13 -962 -9 -956
rect 7 -962 11 -956
rect 15 -962 19 -956
rect -3 -991 1 -982
rect 23 -991 27 -982
rect -27 -994 -12 -991
rect -3 -995 16 -991
rect 23 -995 33 -991
rect -16 -1002 0 -999
rect 7 -1005 11 -995
rect 23 -998 27 -995
rect 15 -1012 19 -1008
rect 19 -1016 25 -1012
rect 11 -1025 33 -1021
rect -13 -1029 -9 -1025
rect -9 -1033 -3 -1029
rect 1 -1033 7 -1029
<< m2contact >>
rect 85 -21 90 -16
rect 118 -29 123 -24
rect 53 -43 58 -38
rect -21 -377 -16 -372
rect -21 -454 -16 -449
rect -21 -559 -16 -554
rect -21 -636 -16 -631
rect -21 -743 -16 -738
rect -21 -820 -16 -815
rect -21 -925 -16 -920
rect -21 -1002 -16 -997
<< metal2 >>
rect 85 -26 89 -21
rect 85 -29 118 -26
rect 85 -43 89 -29
rect 53 -46 89 -43
rect -19 -449 -16 -377
rect -19 -631 -16 -559
rect -19 -815 -16 -743
rect -19 -997 -16 -925
<< labels >>
rlabel space -33 -60 3 19 1 inverter
rlabel space 46 -75 177 26 1 flipflop
rlabel metal1 51 -49 51 -49 1 in_ff
rlabel metal1 51 -40 51 -40 1 clk
rlabel metal1 170 -21 170 -21 1 out_ff
rlabel metal1 -24 -30 -24 -30 1 in_inv
rlabel metal1 -4 -30 -4 -30 1 out_inv
rlabel metal1 -14 9 -14 9 1 vdd
rlabel metal1 238 -66 238 -66 1 gnd
rlabel space 202 -79 293 29 1 xor
rlabel metal1 208 -38 208 -38 1 in2_xor
rlabel metal1 208 -45 208 -45 1 in1_xor
rlabel metal1 284 -45 284 -45 1 out_xor
rlabel metal1 262 -6 262 -6 1 vdd
rlabel space -23 -216 28 -119 1 NAND2
rlabel metal1 4 -129 4 -129 1 vdd
rlabel metal1 -17 -168 -17 -168 1 in1_NAND2
rlabel metal1 -17 -175 -17 -175 1 in2_NAND2
rlabel metal1 4 -206 4 -206 1 gnd
rlabel metal1 15 -168 15 -168 1 out_NAND2
rlabel metal1 54 -168 54 -168 1 in1_NAND3
rlabel metal1 54 -175 54 -175 1 in2_NAND3
rlabel metal1 54 -182 54 -182 1 in3_NAND3
rlabel metal1 76 -129 76 -129 1 vdd
rlabel metal1 76 -223 76 -223 1 gnd
rlabel metal1 98 -175 98 -175 7 out_NAND3
rlabel space 47 -230 104 -117 1 NAND3
rlabel metal1 149 -129 149 -129 1 vdd
rlabel metal1 150 -240 150 -240 1 gnd
rlabel metal1 128 -168 128 -168 1 in1_NAND4
rlabel metal1 128 -175 128 -175 1 in2_NAND4
rlabel metal1 128 -182 128 -182 1 in3_NAND4
rlabel metal1 128 -189 128 -189 1 in4_NAND4
rlabel metal1 184 -175 184 -175 7 out_NAND4
rlabel space 122 -246 190 -120 1 NAND4
rlabel metal1 257 -129 257 -129 1 vdd
rlabel metal1 258 -257 258 -257 1 gnd
rlabel metal1 236 -168 236 -168 1 in1_NAND5
rlabel metal1 236 -175 236 -175 1 in2_NAND5
rlabel metal1 236 -182 236 -182 1 in3_NAND5
rlabel metal1 236 -189 236 -189 1 in4_NAND5
rlabel metal1 236 -196 236 -196 1 in5_NAND5
rlabel metal1 304 -182 304 -182 7 out_NAND5
rlabel metal1 37 -336 37 -336 1 vdd
rlabel metal1 13 -396 13 -396 1 gnd
rlabel metal1 4 -406 4 -406 1 vdd
rlabel metal1 4 -483 4 -483 1 gnd
rlabel metal1 22 -466 22 -466 1 gnd
rlabel metal1 -14 -51 -14 -51 1 gnd
rlabel metal1 22 -648 22 -648 1 gnd
rlabel metal1 4 -665 4 -665 1 gnd
rlabel metal1 4 -588 4 -588 1 vdd
rlabel metal1 13 -578 13 -578 1 gnd
rlabel metal1 37 -518 37 -518 1 vdd
rlabel metal1 37 -702 37 -702 1 vdd
rlabel metal1 13 -762 13 -762 1 gnd
rlabel metal1 4 -772 4 -772 1 vdd
rlabel metal1 4 -849 4 -849 1 gnd
rlabel metal1 22 -832 22 -832 1 gnd
rlabel metal1 22 -1014 22 -1014 1 gnd
rlabel metal1 4 -1031 4 -1031 1 gnd
rlabel metal1 4 -954 4 -954 1 vdd
rlabel metal1 13 -944 13 -944 1 gnd
rlabel metal1 37 -884 37 -884 1 vdd
rlabel metal1 -25 -368 -25 -368 1 a0
rlabel metal2 -18 -380 -18 -380 1 b0
rlabel metal1 59 -375 59 -375 1 p0
rlabel metal1 31 -475 31 -475 1 g0_inv
rlabel metal1 31 -445 31 -445 1 g0
rlabel metal1 -25 -550 -25 -550 1 a1
rlabel metal2 -17 -561 -17 -561 1 b1
rlabel metal1 59 -557 59 -557 1 p1
rlabel metal1 31 -657 31 -657 1 g1_inv
rlabel metal1 31 -627 31 -627 1 g1
rlabel metal1 -25 -734 -25 -734 1 a2
rlabel metal2 -17 -745 -17 -745 1 b2
rlabel metal1 59 -741 59 -741 1 p2
rlabel metal1 31 -811 31 -811 1 g2
rlabel metal1 31 -841 31 -841 1 g2_inv
rlabel metal1 -25 -916 -25 -916 1 a3
rlabel metal2 -17 -927 -17 -927 1 b3
rlabel metal1 59 -923 59 -923 1 p3
rlabel metal1 31 -993 31 -993 1 g3
rlabel metal1 31 -1023 31 -1023 1 g3_inv
<< end >>
