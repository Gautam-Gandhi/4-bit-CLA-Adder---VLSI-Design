magic
tech scmos
timestamp 1731859048
<< nwell >>
rect -26 -25 -2 14
rect 49 -16 172 23
rect 206 -1 246 24
rect 49 -36 85 -16
rect 206 -35 286 -1
rect 246 -40 286 -35
rect -19 -163 17 -124
rect 52 -163 100 -124
rect 126 -163 186 -124
rect 234 -163 306 -124
<< ntransistor >>
rect -15 -45 -13 -35
rect 96 -50 98 -30
rect 108 -50 110 -30
rect 131 -50 133 -30
rect 143 -50 145 -30
rect 159 -36 161 -26
rect 60 -64 62 -54
rect 217 -60 219 -50
rect 257 -60 259 -50
rect 273 -60 275 -50
rect -8 -200 -6 -180
rect 4 -200 6 -180
rect 63 -217 65 -187
rect 75 -217 77 -187
rect 87 -217 89 -187
rect 137 -234 139 -194
rect 149 -234 151 -194
rect 161 -234 163 -194
rect 173 -234 175 -194
rect 245 -251 247 -201
rect 257 -251 259 -201
rect 269 -251 271 -201
rect 281 -251 283 -201
rect 293 -251 295 -201
<< ptransistor >>
rect -15 -19 -13 1
rect 60 -30 62 10
rect 72 -30 74 10
rect 96 -10 98 10
rect 131 -10 133 10
rect 159 -10 161 10
rect 217 -29 219 11
rect 233 -29 235 11
rect 257 -34 259 -14
rect 273 -34 275 -14
rect -8 -157 -6 -137
rect 4 -157 6 -137
rect 63 -157 65 -137
rect 75 -157 77 -137
rect 87 -157 89 -137
rect 137 -157 139 -137
rect 149 -157 151 -137
rect 161 -157 163 -137
rect 173 -157 175 -137
rect 245 -157 247 -137
rect 257 -157 259 -137
rect 269 -157 271 -137
rect 281 -157 283 -137
rect 293 -157 295 -137
<< ndiffusion >>
rect -16 -45 -15 -35
rect -13 -45 -12 -35
rect 95 -50 96 -30
rect 98 -50 108 -30
rect 110 -50 111 -30
rect 130 -50 131 -30
rect 133 -50 143 -30
rect 145 -50 146 -30
rect 158 -36 159 -26
rect 161 -36 162 -26
rect 59 -64 60 -54
rect 62 -64 63 -54
rect 216 -60 217 -50
rect 219 -60 220 -50
rect 256 -60 257 -50
rect 259 -60 260 -50
rect 272 -60 273 -50
rect 275 -60 276 -50
rect -9 -200 -8 -180
rect -6 -200 4 -180
rect 6 -200 7 -180
rect 62 -217 63 -187
rect 65 -217 75 -187
rect 77 -217 87 -187
rect 89 -217 90 -187
rect 136 -234 137 -194
rect 139 -234 149 -194
rect 151 -234 161 -194
rect 163 -234 173 -194
rect 175 -234 176 -194
rect 244 -251 245 -201
rect 247 -251 257 -201
rect 259 -251 269 -201
rect 271 -251 281 -201
rect 283 -251 293 -201
rect 295 -251 296 -201
<< pdiffusion >>
rect -16 -19 -15 1
rect -13 -19 -12 1
rect 59 -30 60 10
rect 62 -30 72 10
rect 74 -30 75 10
rect 95 -10 96 10
rect 98 -10 99 10
rect 130 -10 131 10
rect 133 -10 134 10
rect 158 -10 159 10
rect 161 -10 162 10
rect 216 -29 217 11
rect 219 -29 220 11
rect 232 -29 233 11
rect 235 -29 236 11
rect 256 -34 257 -14
rect 259 -34 260 -14
rect 272 -34 273 -14
rect 275 -34 276 -14
rect -9 -157 -8 -137
rect -6 -157 -5 -137
rect 3 -157 4 -137
rect 6 -157 7 -137
rect 62 -157 63 -137
rect 65 -157 66 -137
rect 74 -157 75 -137
rect 77 -157 78 -137
rect 86 -157 87 -137
rect 89 -157 90 -137
rect 136 -157 137 -137
rect 139 -157 140 -137
rect 148 -157 149 -137
rect 151 -157 152 -137
rect 160 -157 161 -137
rect 163 -157 164 -137
rect 172 -157 173 -137
rect 175 -157 176 -137
rect 244 -157 245 -137
rect 247 -157 248 -137
rect 256 -157 257 -137
rect 259 -157 260 -137
rect 268 -157 269 -137
rect 271 -157 272 -137
rect 280 -157 281 -137
rect 283 -157 284 -137
rect 292 -157 293 -137
rect 295 -157 296 -137
<< ndcontact >>
rect -20 -45 -16 -35
rect -12 -45 -8 -35
rect 91 -50 95 -30
rect 111 -50 115 -30
rect 126 -50 130 -30
rect 146 -50 150 -30
rect 154 -36 158 -26
rect 162 -36 166 -26
rect 55 -64 59 -54
rect 63 -64 67 -54
rect 212 -60 216 -50
rect 220 -60 224 -50
rect 252 -60 256 -50
rect 260 -60 264 -50
rect 268 -60 272 -50
rect 276 -60 280 -50
rect -13 -200 -9 -180
rect 7 -200 11 -180
rect 58 -217 62 -187
rect 90 -217 94 -187
rect 132 -234 136 -194
rect 176 -234 180 -194
rect 240 -251 244 -201
rect 296 -251 300 -201
<< pdcontact >>
rect -20 -19 -16 1
rect -12 -19 -8 1
rect 55 -30 59 10
rect 75 -30 79 10
rect 91 -10 95 10
rect 99 -10 103 10
rect 126 -10 130 10
rect 134 -10 138 10
rect 154 -10 158 10
rect 162 -10 166 10
rect 212 -29 216 11
rect 220 -29 224 11
rect 228 -29 232 11
rect 236 -29 240 11
rect 252 -34 256 -14
rect 260 -34 264 -14
rect 268 -34 272 -14
rect 276 -34 280 -14
rect -13 -157 -9 -137
rect -5 -157 3 -137
rect 7 -157 11 -137
rect 58 -157 62 -137
rect 66 -157 74 -137
rect 78 -157 86 -137
rect 90 -157 94 -137
rect 132 -157 136 -137
rect 140 -157 148 -137
rect 152 -157 160 -137
rect 164 -157 172 -137
rect 176 -157 180 -137
rect 240 -157 244 -137
rect 248 -157 256 -137
rect 260 -157 268 -137
rect 272 -157 280 -137
rect 284 -157 292 -137
rect 296 -157 300 -137
<< psubstratepcontact >>
rect -20 -53 -16 -49
rect -10 -53 -6 -49
rect 154 -44 158 -40
rect 164 -44 168 -40
rect 72 -58 76 -54
rect 87 -58 91 -54
rect 103 -58 107 -54
rect 122 -58 126 -54
rect 138 -58 142 -54
rect 154 -58 158 -54
rect 212 -68 216 -64
rect 220 -68 224 -64
rect 252 -68 256 -64
rect 260 -68 264 -64
rect 268 -68 272 -64
rect 276 -68 280 -64
rect 51 -72 55 -68
rect 62 -72 66 -68
rect 72 -72 76 -68
rect -13 -208 -9 -204
rect -3 -208 1 -204
rect 7 -208 11 -204
rect 58 -225 62 -221
rect 69 -225 73 -221
rect 79 -225 83 -221
rect 90 -225 94 -221
rect 132 -242 136 -238
rect 142 -242 146 -238
rect 154 -242 158 -238
rect 166 -242 170 -238
rect 176 -242 180 -238
rect 240 -259 244 -255
rect 250 -259 254 -255
rect 262 -259 266 -255
rect 274 -259 278 -255
rect 286 -259 290 -255
rect 296 -259 300 -255
<< nsubstratencontact >>
rect 53 16 57 20
rect 65 16 69 20
rect 76 16 80 20
rect 87 16 91 20
rect 101 16 105 20
rect 112 16 116 20
rect 122 16 126 20
rect 136 16 140 20
rect 152 16 156 20
rect 164 16 168 20
rect -22 7 -18 11
rect -10 7 -6 11
rect 252 -8 256 -4
rect 268 -8 272 -4
rect -13 -131 -9 -127
rect -3 -131 1 -127
rect 7 -131 11 -127
rect 58 -131 62 -127
rect 69 -131 73 -127
rect 80 -131 84 -127
rect 90 -131 94 -127
rect 132 -131 136 -127
rect 143 -131 147 -127
rect 154 -131 158 -127
rect 165 -131 169 -127
rect 176 -131 180 -127
rect 240 -131 244 -127
rect 251 -131 255 -127
rect 262 -131 266 -127
rect 273 -131 277 -127
rect 286 -131 290 -127
rect 296 -131 300 -127
<< polysilicon >>
rect 60 10 62 13
rect 72 10 74 13
rect 96 10 98 13
rect 131 10 133 13
rect 159 10 161 13
rect 217 11 219 14
rect 233 11 235 14
rect -15 1 -13 4
rect -15 -35 -13 -19
rect 96 -30 98 -10
rect 108 -30 110 -23
rect 131 -30 133 -10
rect 143 -30 145 -23
rect 159 -26 161 -10
rect -15 -48 -13 -45
rect 60 -54 62 -30
rect 72 -44 74 -30
rect 257 -14 259 -11
rect 273 -14 275 -11
rect 159 -39 161 -36
rect 217 -50 219 -29
rect 233 -40 235 -29
rect 257 -50 259 -34
rect 273 -50 275 -34
rect 96 -53 98 -50
rect 108 -53 110 -50
rect 131 -53 133 -50
rect 143 -53 145 -50
rect 217 -63 219 -60
rect 257 -63 259 -60
rect 273 -63 275 -60
rect 60 -67 62 -64
rect -8 -137 -6 -134
rect 4 -137 6 -134
rect 63 -137 65 -134
rect 75 -137 77 -134
rect 87 -137 89 -134
rect 137 -137 139 -134
rect 149 -137 151 -134
rect 161 -137 163 -134
rect 173 -137 175 -134
rect 245 -137 247 -134
rect 257 -137 259 -134
rect 269 -137 271 -134
rect 281 -137 283 -134
rect 293 -137 295 -134
rect -8 -180 -6 -157
rect 4 -180 6 -157
rect 63 -187 65 -157
rect 75 -187 77 -157
rect 87 -187 89 -157
rect -8 -203 -6 -200
rect 4 -203 6 -200
rect 137 -194 139 -157
rect 149 -194 151 -157
rect 161 -194 163 -157
rect 173 -194 175 -157
rect 63 -220 65 -217
rect 75 -220 77 -217
rect 87 -220 89 -217
rect 245 -201 247 -157
rect 257 -201 259 -157
rect 269 -201 271 -157
rect 281 -201 283 -157
rect 293 -201 295 -157
rect 137 -237 139 -234
rect 149 -237 151 -234
rect 161 -237 163 -234
rect 173 -237 175 -234
rect 245 -254 247 -251
rect 257 -254 259 -251
rect 269 -254 271 -251
rect 281 -254 283 -251
rect 293 -254 295 -251
<< polycontact >>
rect -19 -32 -15 -28
rect 92 -20 96 -16
rect 127 -21 131 -17
rect 104 -27 108 -23
rect 155 -23 159 -19
rect 139 -27 143 -23
rect 56 -51 60 -47
rect 68 -42 72 -38
rect 213 -47 217 -43
rect 229 -40 233 -36
rect 253 -47 257 -43
rect 269 -47 273 -43
rect -12 -170 -8 -166
rect 0 -177 4 -173
rect 59 -170 63 -166
rect 71 -177 75 -173
rect 83 -184 87 -180
rect 133 -170 137 -166
rect 145 -177 149 -173
rect 157 -184 161 -180
rect 169 -191 173 -187
rect 241 -170 245 -166
rect 253 -177 257 -173
rect 265 -184 269 -180
rect 277 -191 281 -187
rect 289 -198 293 -194
<< metal1 >>
rect 49 16 53 20
rect 57 16 65 20
rect 69 16 76 20
rect 80 16 87 20
rect 91 16 101 20
rect 105 16 112 20
rect 116 16 122 20
rect 126 16 136 20
rect 140 16 152 20
rect 156 16 164 20
rect 168 16 172 20
rect 206 17 246 21
rect -26 7 -22 11
rect -18 7 -10 11
rect -6 7 -2 11
rect 55 10 59 16
rect 91 10 95 16
rect 126 10 130 16
rect 154 10 158 16
rect 212 11 216 17
rect 228 11 232 17
rect -20 1 -16 7
rect -12 -28 -8 -19
rect -26 -32 -19 -28
rect -12 -32 -2 -28
rect 90 -20 92 -16
rect 99 -17 103 -10
rect 134 -17 138 -10
rect 99 -20 127 -17
rect 111 -21 127 -20
rect 134 -19 150 -17
rect 162 -19 166 -10
rect 134 -20 155 -19
rect 79 -27 104 -24
rect 111 -30 115 -21
rect 146 -23 155 -20
rect 162 -23 172 -19
rect 123 -27 139 -24
rect 146 -30 150 -23
rect 162 -26 166 -23
rect -12 -35 -8 -32
rect 49 -42 53 -38
rect 58 -42 68 -38
rect -20 -49 -16 -45
rect 75 -47 79 -30
rect -26 -53 -20 -49
rect -16 -53 -10 -49
rect -6 -53 -2 -49
rect 49 -51 56 -47
rect 63 -51 79 -47
rect 221 -36 224 -29
rect 154 -40 158 -36
rect 206 -40 229 -36
rect 158 -44 164 -40
rect 168 -44 172 -40
rect 237 -43 240 -29
rect 63 -54 67 -51
rect 91 -54 95 -50
rect 126 -54 130 -50
rect 154 -54 158 -44
rect 206 -47 213 -43
rect 217 -47 240 -43
rect 243 -43 246 17
rect 256 -8 268 -4
rect 252 -14 256 -8
rect 268 -14 272 -8
rect 260 -43 264 -34
rect 276 -43 280 -34
rect 243 -47 253 -43
rect 260 -47 269 -43
rect 276 -47 286 -43
rect 243 -50 246 -47
rect 260 -50 264 -47
rect 276 -50 280 -47
rect 76 -58 87 -54
rect 91 -58 103 -54
rect 107 -58 122 -54
rect 126 -58 138 -54
rect 142 -58 154 -54
rect 55 -68 59 -64
rect 72 -68 76 -58
rect 224 -53 246 -50
rect 212 -64 216 -60
rect 252 -64 256 -60
rect 268 -64 272 -60
rect 206 -68 212 -64
rect 216 -68 220 -64
rect 224 -68 252 -64
rect 256 -68 260 -64
rect 264 -68 268 -64
rect 272 -68 276 -64
rect 49 -72 51 -68
rect 55 -72 62 -68
rect 66 -72 72 -68
rect -9 -131 -3 -127
rect 1 -131 7 -127
rect -13 -137 -9 -131
rect 7 -137 11 -131
rect 62 -131 69 -127
rect 73 -131 80 -127
rect 84 -131 90 -127
rect 136 -131 143 -127
rect 147 -131 154 -127
rect 158 -131 165 -127
rect 169 -131 176 -127
rect 58 -137 62 -131
rect 80 -137 84 -131
rect 132 -137 136 -131
rect 154 -137 158 -131
rect 176 -137 180 -131
rect 244 -131 251 -127
rect 255 -131 262 -127
rect 266 -131 273 -127
rect 277 -131 286 -127
rect 290 -131 296 -127
rect 240 -137 244 -131
rect 262 -137 266 -131
rect 286 -137 290 -131
rect -3 -166 1 -157
rect 68 -166 72 -157
rect 90 -166 94 -157
rect 142 -160 146 -157
rect 166 -160 170 -157
rect 142 -163 170 -160
rect 250 -160 254 -157
rect 274 -160 278 -157
rect 296 -160 300 -157
rect 250 -163 300 -160
rect -19 -170 -12 -166
rect -3 -170 17 -166
rect 52 -170 59 -166
rect 68 -170 94 -166
rect 126 -170 133 -166
rect -19 -177 0 -173
rect 7 -180 11 -170
rect 90 -173 94 -170
rect 166 -173 170 -163
rect 234 -170 241 -166
rect 52 -177 71 -173
rect 90 -177 100 -173
rect 126 -177 145 -173
rect 166 -177 186 -173
rect 234 -177 253 -173
rect 52 -184 83 -180
rect 90 -187 94 -177
rect 126 -184 157 -180
rect -13 -204 -9 -200
rect -9 -208 -3 -204
rect 1 -208 7 -204
rect 126 -191 169 -187
rect 176 -194 180 -177
rect 296 -180 300 -163
rect 234 -184 265 -180
rect 296 -184 306 -180
rect 234 -191 277 -187
rect 58 -221 62 -217
rect 62 -225 69 -221
rect 73 -225 79 -221
rect 83 -225 90 -221
rect 234 -198 289 -194
rect 296 -201 300 -184
rect 132 -238 136 -234
rect 136 -242 142 -238
rect 146 -242 154 -238
rect 158 -242 166 -238
rect 170 -242 176 -238
rect 240 -255 244 -251
rect 244 -259 250 -255
rect 254 -259 262 -255
rect 266 -259 274 -255
rect 278 -259 286 -255
rect 290 -259 296 -255
<< m2contact >>
rect 85 -21 90 -16
rect 118 -29 123 -24
rect 53 -43 58 -38
<< metal2 >>
rect 85 -26 89 -21
rect 85 -29 118 -26
rect 85 -43 89 -29
rect 53 -46 89 -43
<< labels >>
rlabel space -33 -60 3 19 1 inverter
rlabel space 46 -75 177 26 1 flipflop
rlabel metal1 51 -49 51 -49 1 in_ff
rlabel metal1 51 -40 51 -40 1 clk
rlabel metal1 170 -21 170 -21 1 out_ff
rlabel metal1 -24 -30 -24 -30 1 in_inv
rlabel metal1 -4 -30 -4 -30 1 out_inv
rlabel metal1 -14 9 -14 9 1 vdd
rlabel metal1 -13 -51 -13 -51 1 gnd
rlabel metal1 238 -66 238 -66 1 gnd
rlabel space 202 -79 293 29 1 xor
rlabel metal1 208 -38 208 -38 1 in2_xor
rlabel metal1 208 -45 208 -45 1 in1_xor
rlabel metal1 284 -45 284 -45 1 out_xor
rlabel metal1 262 -6 262 -6 1 vdd
rlabel space -23 -216 28 -119 1 NAND2
rlabel metal1 4 -129 4 -129 1 vdd
rlabel metal1 -17 -168 -17 -168 1 in1_NAND2
rlabel metal1 -17 -175 -17 -175 1 in2_NAND2
rlabel metal1 4 -206 4 -206 1 gnd
rlabel metal1 15 -168 15 -168 1 out_NAND2
rlabel metal1 54 -168 54 -168 1 in1_NAND3
rlabel metal1 54 -175 54 -175 1 in2_NAND3
rlabel metal1 54 -182 54 -182 1 in3_NAND3
rlabel metal1 76 -129 76 -129 1 vdd
rlabel metal1 76 -223 76 -223 1 gnd
rlabel metal1 98 -175 98 -175 7 out_NAND3
rlabel space 47 -230 104 -117 1 NAND3
rlabel metal1 149 -129 149 -129 1 vdd
rlabel metal1 150 -240 150 -240 1 gnd
rlabel metal1 128 -168 128 -168 1 in1_NAND4
rlabel metal1 128 -175 128 -175 1 in2_NAND4
rlabel metal1 128 -182 128 -182 1 in3_NAND4
rlabel metal1 128 -189 128 -189 1 in4_NAND4
rlabel metal1 184 -175 184 -175 7 out_NAND4
rlabel space 122 -246 190 -120 1 NAND4
rlabel metal1 257 -129 257 -129 1 vdd
rlabel metal1 258 -257 258 -257 1 gnd
rlabel metal1 236 -168 236 -168 1 in1_NAND5
rlabel metal1 236 -175 236 -175 1 in2_NAND5
rlabel metal1 236 -182 236 -182 1 in3_NAND5
rlabel metal1 236 -189 236 -189 1 in4_NAND5
rlabel metal1 236 -196 236 -196 1 in5_NAND5
rlabel metal1 304 -182 304 -182 7 out_NAND5
<< end >>
