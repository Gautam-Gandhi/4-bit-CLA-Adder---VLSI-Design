* SPICE3 file created from NAND3.ext - technology: scmos

.option scale=90n

M1000 out_xor a_21_n168# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1001 a_n26_n137# in1_xor gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1002 a_62_n30# in_ff w_49_n36# w_49_n36# pfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1003 in1_xor in2_xor a_n26_n137# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1004 a_62_n64# clk a_62_n30# w_49_n36# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1005 a_98_n10# clk w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1006 out_inv in_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1007 a_157_n202# in1_NAND3 gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1008 out_xor a_21_n168# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1009 out_NAND3 in1_NAND3 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1010 a_86_n185# in1_NAND2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1011 out_inv in_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1012 out_ff a_133_n10# a_51_n72# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1013 a_21_n168# a_n26_n137# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 a_169_n202# in2_NAND3 a_157_n202# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1015 in2_xor in1_xor a_n26_n137# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1016 a_133_n50# a_98_n10# a_51_n72# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1017 vdd in2_NAND3 out_NAND3 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1018 a_98_n50# clk a_51_n72# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1019 a_98_n10# a_62_n64# a_98_n50# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1020 out_NAND2 in2_NAND2 a_86_n185# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1021 a_62_n64# in_ff a_51_n72# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1022 out_NAND2 in1_NAND2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1023 a_133_n10# a_98_n10# w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1024 out_NAND3 in3_NAND3 a_169_n202# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1025 a_133_n10# clk a_133_n50# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1026 out_ff a_133_n10# w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1027 out_NAND3 in3_NAND3 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1028 vdd in2_NAND2 out_NAND2 vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1029 a_21_n168# a_n26_n137# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
C0 a_98_n10# a_62_n64# 0.163856f
C1 in_inv out_inv 0.059344f
C2 vdd out_NAND3 0.662121f
C3 w_49_n36# clk 0.069031f
C4 clk a_133_n50# 1.7e-19
C5 a_133_n10# a_51_n72# 0.304049f
C6 vdd in2_xor 0.02552f
C7 in1_xor in2_xor 0.424419f
C8 out_inv gnd 0.123737f
C9 gnd in1_NAND3 0.001614f
C10 gnd a_157_n202# 1.36e-19
C11 w_49_n36# a_98_n10# 0.272577f
C12 a_21_n168# out_xor 0.059344f
C13 vdd a_n26_n137# 0.317981f
C14 in1_xor a_n26_n137# 1.51355f
C15 gnd in2_NAND3 8.87e-19
C16 a_133_n10# out_ff 0.059344f
C17 gnd a_169_n202# 1.36e-19
C18 in_ff clk 0.125563f
C19 w_49_n36# a_133_n10# 0.248779f
C20 in1_NAND3 in2_NAND3 0.173673f
C21 vdd a_21_n168# 0.467651f
C22 in2_xor a_n26_n137# 0.90085f
C23 gnd in3_NAND3 0.0559f
C24 in1_NAND3 in3_NAND3 0.007681f
C25 in1_NAND2 out_NAND2 0.036296f
C26 vdd in1_NAND2 0.020614f
C27 a_157_n202# in3_NAND3 2.83e-19
C28 gnd out_xor 0.103118f
C29 clk a_98_n10# 0.33274f
C30 vdd in_inv 0.020614f
C31 in2_NAND3 in3_NAND3 0.339028f
C32 in2_NAND2 out_NAND2 0.163729f
C33 vdd in2_NAND2 0.020473f
C34 a_62_n64# a_51_n72# 0.260028f
C35 a_n26_n137# a_21_n168# 0.059344f
C36 a_51_n72# a_98_n50# 1.36e-19
C37 gnd out_NAND2 2.27e-20
C38 a_169_n202# in3_NAND3 1.7e-19
C39 gnd in1_xor 0.056598f
C40 w_49_n36# a_62_n30# 6.79e-20
C41 clk a_133_n10# 0.163856f
C42 vdd out_inv 0.22794f
C43 out_ff a_51_n72# 0.123737f
C44 a_62_n64# a_98_n50# 1.7e-19
C45 vdd in1_NAND3 0.020614f
C46 a_51_n72# a_133_n50# 1.36e-19
C47 gnd out_NAND3 2.27e-20
C48 w_49_n36# a_62_n64# 0.020872f
C49 a_98_n10# a_133_n10# 0.044023f
C50 in1_NAND3 out_NAND3 0.036296f
C51 vdd in2_NAND3 0.020472f
C52 gnd a_n26_n137# 0.180335f
C53 w_49_n36# out_ff 0.22794f
C54 in2_NAND3 out_NAND3 0.106322f
C55 vdd in3_NAND3 0.020472f
C56 in_ff a_51_n72# 0.056598f
C57 gnd a_21_n168# 0.262811f
C58 in_ff a_62_n64# 0.057163f
C59 in3_NAND3 out_NAND3 0.069367f
C60 vdd out_xor 0.214182f
C61 in1_NAND2 in2_NAND2 0.174076f
C62 clk a_51_n72# 0.059299f
C63 gnd in1_NAND2 0.001614f
C64 a_86_n185# in2_NAND2 1.7e-19
C65 a_86_n185# gnd 1.36e-19
C66 clk a_62_n64# 0.341152f
C67 vdd out_NAND2 0.448048f
C68 w_49_n36# in_ff 0.020473f
C69 vdd in1_xor 0.024924f
C70 clk a_98_n50# 5.16e-20
C71 a_98_n10# a_51_n72# 0.042875f
C72 in_inv gnd 0.056598f
C73 gnd in2_NAND2 0.0559f
