* SPICE3 file created from cla.ext - technology: scmos

.option scale=90n

M1000 c4 g3_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1001 a_100_n781# c0 a_88_n781# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1002 a_110_n1392# a_116_n1412# a_110_n1435# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1003 vdd a_94_n825# c3 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1004 out_NAND3 in1_NAND3 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1005 g1 g1_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1006 a_118_n1118# c0 a_106_n1118# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1007 p2 a_34_n808# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1008 g1_inv a1 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1009 g1_inv b1 a_n6_n659# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1010 c2 a_82_n504# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1011 a_88_n704# p0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1012 p2 c2 a_151_n725# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1013 out_xor a_259_n60# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1014 vdd p2 a_100_n1287# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1015 a_100_n1347# g1 gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1016 a_94_n825# p2 a_106_n885# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1017 a_82_n504# p1 a_94_n564# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1018 vdd b2 g2_inv vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1019 s3 a_268_n808# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1020 a_62_n30# in_ff w_49_n36# w_49_n36# pfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1021 in1_xor in2_xor a_212_n29# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1022 out_NAND4 in4_NAND4 a_163_n234# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1023 p1 a_34_n572# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1024 a_158_n845# a_88_n704# gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1025 a_100_n1287# p3 a_112_n1347# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1026 a_77_n217# in2_NAND3 a_65_n217# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1027 a_110_n1435# p3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1028 a_n13_n541# b1 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1029 g2 g2_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1030 vdd in2_NAND5 out_NAND5 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1031 c0 p0 a_150_n403# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1032 g3_inv b3 a_n6_n1276# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1033 a_100_n1287# g1 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1034 a_62_n64# clk a_62_n30# w_49_n36# pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1035 c1 p1 a_169_n498# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1036 a_136_n564# a_82_n504# gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1037 vdd in2_NAND4 out_NAND4 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1038 a_82_n1024# p3 a_118_n1118# Gnd nfet w=50 l=2
+  ad=0.25n pd=0.11m as=0.25n ps=60u
M1039 s1 a_216_n473# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1040 vdd a_90_n1164# c4 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1041 vdd p1 a_90_n1164# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1042 a_100_n1287# p3 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1043 vdd in2_NAND3 out_NAND3 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1044 a_216_n473# a_169_n498# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1045 s3 a_268_n808# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1046 a_169_n498# c1 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1047 vdd a_82_n608# c2 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1048 a2 b2 a_n13_n777# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1049 a_98_n10# clk w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1050 vdd p1 a_88_n704# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1051 a_82_n1024# p2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1052 a_139_n234# in1_NAND4 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1053 a_34_n383# a_n13_n352# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1054 out_inv in_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1055 p3 c3 a_221_n777# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1056 a_259_n60# a_212_n29# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1057 vdd b1 g1_inv vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1058 a_170_n845# a_94_n825# a_158_n845# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1059 out_NAND3 in3_NAND3 a_77_n217# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1060 a_108_n400# a_73_n357# gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1061 c4 a_82_n1024# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1062 in2_xor in1_xor a_212_n29# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1063 a_90_n1164# p2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1064 a_88_n704# p2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1065 a_n6_n1276# a3 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1066 g1 g1_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1067 out_NAND5 in3_NAND5 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1068 c4 g3_inv a_197_n1258# Gnd nfet w=50 l=2
+  ad=0.25n pd=0.11m as=0.25n ps=60u
M1069 p3 a_34_n1189# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1070 a_n13_n1158# b3 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1071 c4 a_100_n1287# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1072 a_90_n1164# p3 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1073 a_148_n564# a_82_n608# a_136_n564# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1074 a0 b0 a_n13_n352# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1075 a_n13_n777# b2 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1076 a_73_n400# p0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1077 a_34_n1189# a_n13_n1158# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1078 vdd b3 g3_inv vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1079 out_NAND3 in3_NAND3 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1080 vdd p1 a_82_n1024# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1081 a_283_n251# in4_NAND5 a_271_n251# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1082 p0 a_34_n383# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1083 c2 g1_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1084 b2 a2 a_n13_n777# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1085 out_xor a_259_n60# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1086 a_151_n234# in2_NAND4 a_139_n234# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1087 g3 g3_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1088 a_n6_n470# a0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1089 a_n6_n200# in1_NAND2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1090 a_102_n1241# p1 a_90_n1241# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1091 a_94_n825# p1 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1092 c3 a_94_n929# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1093 c2 p2 a_151_n725# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1094 a_82_n504# c0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1095 c1 g0_inv a_108_n400# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1096 vdd a_116_n1412# a_110_n1392# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1097 vdd c0 a_88_n704# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1098 vdd a_110_n1392# c4 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1099 vdd g0 a_90_n1164# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1100 a_94_n929# p2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1101 c1 a_73_n357# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1102 a_82_n608# g0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1103 a_173_n1258# a_90_n1164# a_161_n1258# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1104 g2 g2_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1105 a_82_n1024# p0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1106 a_112_n781# p0 a_100_n781# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1107 c2 g1_inv a_148_n564# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=0.15n ps=40u
M1108 a_34_n383# a_n13_n352# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1109 a_198_n700# a_151_n725# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1110 g3_inv a3 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1111 out_inv in_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1112 a_73_n357# c0 a_73_n400# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1113 a_90_n1241# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1114 a_82_n1118# p2 gnd Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=0.11m
M1115 a_94_n972# p2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1116 out_ff a_133_n10# a_51_n72# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1117 p0 c0 a_150_n403# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1118 a_82_n651# g0 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1119 a_247_n251# in1_NAND5 gnd Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=0.11m
M1120 b0 a0 a_n13_n352# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1121 a_110_n1392# p3 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1122 b3 a3 a_n13_n1158# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1123 a_94_n885# p1 gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1124 a_n6_n895# a2 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1125 out_NAND5 in5_NAND5 a_283_n251# Gnd nfet w=50 l=2
+  ad=0.25n pd=0.11m as=0.25n ps=60u
M1126 a_34_n572# a_n13_n541# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1127 a_82_n564# c0 gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1128 a_114_n1241# p3 a_102_n1241# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1129 a_73_n357# p0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1130 a_161_n1258# a_82_n1024# gnd Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=0.11m
M1131 out_NAND4 in3_NAND4 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1132 a_268_n808# a_221_n777# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1133 s1 a_216_n473# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1134 vdd p0 a_82_n504# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1135 vdd g2_inv c3 vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1136 a_259_n60# a_212_n29# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1137 a_197_n378# a_150_n403# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1138 g0 g0_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1139 g0_inv b0 a_n6_n470# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1140 a_185_n1258# a_100_n1287# a_173_n1258# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1141 a_212_n29# in1_xor gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1142 out_NAND2 in1_NAND2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1143 out_NAND2 in2_NAND2 a_n6_n200# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1144 g0_inv a0 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1145 vdd c0 a_82_n1024# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1146 a_198_n700# a_151_n725# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1147 a_34_n808# a_n13_n777# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1148 a_133_n50# a_98_n10# a_51_n72# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1149 vdd g0_inv c1 vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1150 vdd p1 a_82_n608# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1151 p0 a_34_n383# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1152 a_98_n50# clk a_51_n72# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1153 a_98_n10# a_62_n64# a_98_n50# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1154 a1 b1 a_n13_n541# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1155 s2 a_198_n700# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1156 a_94_n1118# p1 a_82_n1118# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1157 a_182_n845# a_94_n929# a_170_n845# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1158 a_88_n704# p1 a_112_n781# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1159 vdd g0 a_94_n825# vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1160 p1 c1 a_169_n498# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1161 a_151_n725# c2 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1162 a_n13_n352# b0 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1163 p1 a_34_n572# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1164 a_62_n64# in_ff a_51_n72# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1165 a_259_n251# in2_NAND5 a_247_n251# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1166 a_216_n473# a_169_n498# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1167 a_82_n608# p1 a_82_n651# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1168 a_90_n1164# g0 a_114_n1241# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1169 vdd in4_NAND5 out_NAND5 vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=30u
M1170 vdd g1 a_94_n929# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1171 a_94_n564# p0 a_82_n564# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1172 a_268_n808# a_221_n777# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1173 a_n6_n659# a1 gnd Gnd nfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1174 a_133_n10# a_98_n10# w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1175 vdd c0 a_73_n357# vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1176 a_133_n10# clk a_133_n50# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1177 vdd in4_NAND4 out_NAND4 vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1178 a_197_n378# a_150_n403# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1179 a_88_n781# p2 gnd Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=90u
M1180 g2_inv b2 a_n6_n895# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1181 c3 a_88_n704# vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1182 a_197_n1258# a_110_n1392# a_185_n1258# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1183 g3 g3_inv gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1184 g2_inv a2 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1185 c3 p3 a_221_n777# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1186 s0 a_197_n378# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1187 a_94_n929# g1 a_94_n972# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1188 a_82_n1024# p3 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1189 a_106_n1118# p0 a_94_n1118# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1190 a_34_n808# a_n13_n777# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1191 a_150_n403# p0 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1192 a_106_n885# g0 a_94_n885# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1193 p2 a_34_n808# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1194 out_ff a_133_n10# w_49_n36# w_49_n36# pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1195 s2 a_198_n700# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1196 a_163_n234# in3_NAND4 a_151_n234# Gnd nfet w=40 l=2
+  ad=0.2n pd=50u as=0.2n ps=50u
M1197 a_34_n572# a_n13_n541# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1198 a_65_n217# in1_NAND3 gnd Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=70u
M1199 vdd b0 g0_inv vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1200 c3 g2_inv a_182_n845# Gnd nfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=50u
M1201 vdd in2_NAND2 out_NAND2 vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1202 a_94_n825# p2 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1203 b1 a1 a_n13_n541# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1204 a_82_n504# p1 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1205 a_112_n1347# p2 a_100_n1347# Gnd nfet w=30 l=2
+  ad=0.15n pd=40u as=0.15n ps=40u
M1206 p3 a_34_n1189# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1207 a3 b3 a_n13_n1158# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1208 out_NAND5 in1_NAND5 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1209 a_271_n251# in3_NAND5 a_259_n251# Gnd nfet w=50 l=2
+  ad=0.25n pd=60u as=0.25n ps=60u
M1210 out_NAND5 in5_NAND5 vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=30u
M1211 g0 g0_inv vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1212 out_NAND4 in1_NAND4 vdd vdd pfet w=20 l=2
+  ad=100p pd=30u as=100p ps=50u
M1213 s0 a_197_n378# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1214 a_34_n1189# a_n13_n1158# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1215 a_221_n777# p3 gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
C0 w_49_n36# a_62_n30# 6.79e-20
C1 vdd out_inv 0.214194f
C2 c0 g1_inv 0.004427f
C3 c1 p1 0.590519f
C4 s2 gnd 0.103118f
C5 in5_NAND5 a_283_n251# 1.7e-19
C6 b0 a_n13_n352# 1.51355f
C7 gnd a_139_n234# 1.36e-19
C8 in1_NAND5 in5_NAND5 0.007681f
C9 in2_NAND5 in4_NAND5 0.007278f
C10 g1_inv gnd 0.825349f
C11 a_106_n1118# p3 2.83e-19
C12 a_94_n564# gnd 1.36e-19
C13 a_110_n1392# p3 0.036296f
C14 a_100_n1347# gnd 1.36e-19
C15 g0 vdd 0.30663f
C16 in2_NAND3 out_NAND3 0.106322f
C17 out_xor gnd 0.103118f
C18 gnd out_inv 0.103118f
C19 vdd a_221_n777# 0.31023f
C20 a_90_n1164# a_82_n1024# 0.311133f
C21 g1 p1 0.292837f
C22 a3 a_n13_n1158# 0.90085f
C23 a_34_n383# vdd 0.467651f
C24 a_90_n1164# c4 0.00699f
C25 a_100_n1287# g3_inv 0.00908f
C26 p1 a_116_n1412# 0.26712f
C27 g2_inv a_158_n845# 2.83e-19
C28 vdd b0 0.067865f
C29 gnd a_94_n885# 1.36e-19
C30 a_221_n777# a_268_n808# 0.059344f
C31 in2_NAND5 vdd 0.020472f
C32 in_ff a_62_n64# 0.057163f
C33 a_173_n1258# gnd 1.36e-19
C34 c0 g0 0.049817f
C35 g0 gnd 0.12832f
C36 a_198_n700# vdd 0.467651f
C37 a_94_n929# g2_inv 3.23943f
C38 b2 a_n6_n895# 1.7e-19
C39 gnd a_221_n777# 0.180335f
C40 a_82_n608# vdd 0.46852f
C41 in_ff clk 0.125563f
C42 in1_NAND3 in3_NAND3 0.007681f
C43 p0 c1 0.00227f
C44 a_n13_n1158# vdd 0.31023f
C45 a_34_n383# gnd 0.262811f
C46 a_100_n1287# p2 0.106322f
C47 c3 a_94_n825# 0.00699f
C48 a_88_n781# gnd 1.36e-19
C49 a_n6_n200# gnd 1.36e-19
C50 p1 a_82_n1024# 0.00699f
C51 a_98_n50# a_51_n72# 1.36e-19
C52 in2_NAND4 vdd 0.020472f
C53 a_133_n10# a_51_n72# 0.304049f
C54 g0 g1_inv 0.001428f
C55 a_34_n1189# g1 7.95e-20
C56 in2_NAND5 gnd 8.87e-19
C57 gnd b0 0.114196f
C58 in4_NAND5 out_NAND5 0.007111f
C59 vdd m2_37_n508# 1.53e-19
C60 a_259_n60# vdd 0.467651f
C61 vdd in_inv 0.020614f
C62 p2 a_34_n808# 0.059949f
C63 g1 g2_inv 0.010922f
C64 a_198_n700# gnd 0.262811f
C65 in5_NAND5 a_271_n251# 2.83e-19
C66 b0 a0 0.626439f
C67 p1 a_94_n825# 0.036296f
C68 in1_NAND5 in4_NAND5 0.007278f
C69 gnd a_77_n217# 1.36e-19
C70 in2_NAND5 in3_NAND5 0.338625f
C71 a_82_n608# gnd 9.1e-19
C72 a_94_n1118# p3 2.83e-19
C73 g1 p0 0.12482f
C74 a_n13_n1158# gnd 0.180335f
C75 a_34_n1189# a_116_n1412# 1.09e-20
C76 g1 p3 0.106409f
C77 a_82_n564# gnd 1.36e-19
C78 in4_NAND4 a_163_n234# 1.7e-19
C79 g2_inv a_116_n1412# 0.001471f
C80 in2_NAND4 gnd 8.87e-19
C81 a_151_n725# p2 0.90085f
C82 a_198_n700# s2 0.059344f
C83 a_100_n1287# vdd 0.693459f
C84 a_82_n608# g1_inv 1.32187f
C85 p3 a_116_n1412# 0.346186f
C86 in1_NAND3 out_NAND3 0.036296f
C87 a_259_n60# gnd 0.262811f
C88 gnd in_inv 0.056598f
C89 a_197_n378# vdd 0.467651f
C90 vdd a_34_n808# 0.467651f
C91 out_NAND5 vdd 1.35816f
C92 a_90_n1164# g3_inv 0.007681f
C93 p0 a_82_n1024# 0.007111f
C94 g2_inv g2 0.059062f
C95 p3 a_82_n1024# 0.167001f
C96 gnd a_n6_n895# 1.36e-19
C97 in1_NAND5 vdd 0.020614f
C98 a_100_n1287# gnd 0.012692f
C99 a_110_n1392# a_116_n1412# 0.163729f
C100 a_108_n400# gnd 1.36e-19
C101 a_151_n725# vdd 0.622545f
C102 a_94_n825# g2_inv 0.007681f
C103 a_82_n504# vdd 0.682855f
C104 in1_NAND3 in2_NAND3 0.173673f
C105 p0 g0_inv 0.004837f
C106 out_ff a_51_n72# 0.123737f
C107 a_197_n378# gnd 0.262811f
C108 a_34_n572# vdd 0.467651f
C109 a_90_n1164# p2 0.001572f
C110 a2 g2_inv 0.036296f
C111 out_NAND5 gnd 2.27e-20
C112 a_34_n808# gnd 0.262811f
C113 a_259_n60# out_xor 0.059344f
C114 a_110_n1392# a_82_n1024# 0.007278f
C115 in1_NAND4 vdd 0.020614f
C116 a_133_n10# out_ff 0.059344f
C117 in_inv out_inv 0.059344f
C118 a_98_n10# a_51_n72# 0.042875f
C119 g0 a_82_n608# 0.036296f
C120 gnd a_283_n251# 1.36e-19
C121 in3_NAND5 out_NAND5 0.007111f
C122 in1_NAND5 gnd 0.001614f
C123 g3_inv p1 8.39e-22
C124 a_133_n50# clk 1.7e-19
C125 a_110_n1392# c4 0.007111f
C126 a_212_n29# vdd 0.31023f
C127 a_98_n10# a_133_n10# 0.044023f
C128 g3_inv a_185_n1258# 2.83e-19
C129 a_102_n1241# gnd 1.36e-19
C130 vdd in2_xor 0.02552f
C131 g1 a_94_n929# 0.163729f
C132 c0 a_82_n504# 0.036296f
C133 a_151_n725# gnd 0.180335f
C134 in5_NAND5 a_259_n251# 2.83e-19
C135 in1_NAND5 in3_NAND5 0.007278f
C136 p1 a_112_n781# 1.7e-19
C137 gnd a_65_n217# 1.36e-19
C138 a_82_n504# gnd 0.001637f
C139 a_82_n1118# p3 2.83e-19
C140 a_34_n572# gnd 0.261924f
C141 in4_NAND4 a_151_n234# 2.83e-19
C142 g0 m2_37_n508# 0.021002f
C143 in1_NAND4 gnd 0.001614f
C144 a_90_n1164# vdd 1.041242f
C145 p2 p1 0.922401f
C146 a_82_n504# g1_inv 0.007681f
C147 a_212_n29# gnd 0.180335f
C148 a_169_n498# p1 0.90085f
C149 a_150_n403# vdd 0.310109f
C150 vdd c3 1.04629f
C151 out_NAND4 vdd 1.02077f
C152 g1 a_116_n1412# 0.165053f
C153 in4_NAND4 vdd 0.020473f
C154 gnd a_182_n845# 1.36e-19
C155 vdd m2_67_n574# 2.15e-19
C156 a_118_n1118# p3 1.7e-19
C157 a_90_n1164# gnd 9.1e-19
C158 c0 a_73_n400# 1.7e-19
C159 g0_inv c1 0.163246f
C160 a_73_n400# gnd 1.36e-19
C161 a_94_n825# a_94_n929# 1.17713f
C162 g3_inv p3 5.94e-19
C163 a_112_n1347# gnd 1.36e-19
C164 p1 vdd 0.439582f
C165 w_49_n36# in_ff 0.020473f
C166 p0 a_73_n357# 0.039474f
C167 a_150_n403# c0 1.58815f
C168 a_62_n64# a_51_n72# 0.260028f
C169 a_150_n403# gnd 0.228446f
C170 b2 g2_inv 0.153419f
C171 out_NAND4 gnd 2.27e-20
C172 c3 gnd 2.27e-20
C173 g0 a_102_n1241# 2.83e-19
C174 a_98_n50# a_62_n64# 1.7e-19
C175 in3_NAND3 vdd 0.020472f
C176 clk a_51_n72# 0.059299f
C177 c0 m2_67_n574# 0.01305f
C178 p2 g2_inv 0.001371f
C179 a_88_n704# c3 0.001572f
C180 a2 a_n13_n777# 0.90085f
C181 in2_NAND5 out_NAND5 0.00699f
C182 gnd a_271_n251# 1.36e-19
C183 m2_67_n574# gnd 2.88e-19
C184 in4_NAND4 gnd 0.0559f
C185 a_98_n50# clk 5.16e-20
C186 p2 p0 0.09361f
C187 a_110_n1392# g3_inv 1.24759f
C188 clk a_133_n10# 0.163856f
C189 vdd in1_xor 0.024924f
C190 c0 p1 0.951731f
C191 p2 p3 0.546269f
C192 a_82_n651# gnd 1.36e-19
C193 in5_NAND5 a_247_n251# 2.83e-19
C194 p1 a_100_n781# 2.83e-19
C195 in1_NAND5 in2_NAND5 0.173673f
C196 p1 gnd 0.944202f
C197 a_116_n1412# g2 0.007609f
C198 a_185_n1258# gnd 1.36e-19
C199 p2 c2 0.442092f
C200 in4_NAND4 a_139_n234# 2.83e-19
C201 p1 a_88_n704# 0.070534f
C202 a1 a_n13_n541# 0.90085f
C203 in3_NAND3 gnd 0.0559f
C204 a_151_n725# a_198_n700# 0.059344f
C205 a_n6_n659# b1 1.7e-19
C206 a_34_n1189# vdd 0.467651f
C207 p1 g1_inv 0.004254f
C208 a_82_n504# a_82_n608# 0.737259f
C209 a_169_n498# c2 0.247428f
C210 s0 vdd 0.214182f
C211 in2_NAND2 out_NAND2 0.163729f
C212 gnd in1_xor 0.056598f
C213 vdd g2_inv 0.489553f
C214 g3_inv b3 0.153419f
C215 c4 a_82_n1024# 0.001572f
C216 a_94_n564# p1 1.7e-19
C217 a_216_n473# s1 0.059344f
C218 p0 vdd 0.367036f
C219 a_90_n1164# g0 0.071017f
C220 vdd p3 0.361724f
C221 out_NAND3 vdd 0.662121f
C222 g3_inv g3 0.135151f
C223 in3_NAND4 vdd 0.020472f
C224 gnd a_170_n845# 1.36e-19
C225 c2 vdd 0.687693f
C226 a_90_n1241# gnd 1.36e-19
C227 a_34_n1189# gnd 0.262811f
C228 in1_NAND4 in2_NAND4 0.173673f
C229 a_73_n357# c1 0.036296f
C230 c0 g2_inv 0.007772f
C231 s0 gnd 0.103118f
C232 c3 a_221_n777# 0.90085f
C233 g2_inv gnd 1.103215f
C234 p0 c0 1.64773f
C235 a_110_n1392# vdd 0.468954f
C236 a3 b3 0.626439f
C237 a_n6_n1276# b3 1.7e-19
C238 c0 p3 0.580912f
C239 g0 m2_67_n574# 0.008155f
C240 p0 gnd 0.164553f
C241 g1 a_94_n972# 1.7e-19
C242 a_88_n704# g2_inv 0.007681f
C243 p3 gnd 0.766349f
C244 out_NAND3 gnd 2.27e-20
C245 a_212_n29# a_259_n60# 0.059344f
C246 in2_NAND3 vdd 0.020472f
C247 a_98_n10# a_62_n64# 0.163856f
C248 p0 a_88_n704# 0.010538f
C249 g0 p1 0.529842f
C250 p2 a_94_n929# 0.036296f
C251 b2 a_n13_n777# 1.51355f
C252 g3_inv g1 3.56e-19
C253 in1_NAND5 out_NAND5 0.001572f
C254 gnd a_259_n251# 1.36e-19
C255 in3_NAND4 gnd 8.87e-19
C256 c2 gnd 0.437582f
C257 clk a_98_n10# 0.33274f
C258 a_106_n1118# gnd 1.36e-19
C259 p0 g1_inv 9.7e-19
C260 c1 a_169_n498# 1.51355f
C261 a_n6_n659# gnd 1.36e-19
C262 p1 a_88_n781# 2.83e-19
C263 a_n6_n470# gnd 1.36e-19
C264 a_110_n1392# gnd 9.1e-19
C265 g3_inv a_116_n1412# 0.001561f
C266 vdd b3 0.067865f
C267 b1 a_n13_n541# 1.51355f
C268 g1_inv c2 0.068884f
C269 p3 a_100_n1347# 2.83e-19
C270 a_116_n1412# a_110_n1435# 1.7e-19
C271 in2_NAND4 out_NAND4 0.00699f
C272 in2_NAND3 gnd 8.87e-19
C273 g1 p2 0.58148f
C274 g3 vdd 0.227819f
C275 p1 a_82_n608# 0.163729f
C276 c1 vdd 0.472851f
C277 in1_NAND2 out_NAND2 0.036296f
C278 in2_NAND4 in4_NAND4 0.007681f
C279 vdd a_94_n929# 0.46852f
C280 g3_inv a_82_n1024# 0.007681f
C281 a_82_n564# p1 2.83e-19
C282 a_90_n1164# a_100_n1287# 1.27335f
C283 in3_NAND3 a_77_n217# 1.7e-19
C284 a_90_n1241# g0 6.13e-20
C285 vdd a_n13_n777# 0.31023f
C286 gnd b3 0.114196f
C287 out_NAND2 vdd 0.448048f
C288 g3_inv a_197_n1258# 1.7e-19
C289 g3_inv c4 0.071424f
C290 a_114_n1241# gnd 1.36e-19
C291 g0 g2_inv 5.95e-19
C292 gnd a_158_n845# 1.36e-19
C293 g3 gnd 0.123737f
C294 a_n13_n541# vdd 0.31023f
C295 p0 g0 0.441021f
C296 a_73_n357# g0_inv 0.272103f
C297 c0 c1 0.00147f
C298 g0 p3 0.215667f
C299 c1 gnd 0.053259f
C300 p2 a_82_n1024# 0.001572f
C301 g1 vdd 0.27766f
C302 p3 a_221_n777# 1.51355f
C303 a_94_n929# gnd 9.1e-19
C304 s1 vdd 0.214182f
C305 p0 a_34_n383# 0.059344f
C306 a_150_n403# a_197_n378# 0.059344f
C307 a_88_n704# a_94_n929# 0.007278f
C308 a_n13_n777# gnd 0.180335f
C309 out_NAND2 gnd 2.27e-20
C310 a_212_n29# in2_xor 0.90085f
C311 in1_NAND3 vdd 0.020614f
C312 vdd a_116_n1412# 0.020502f
C313 clk a_62_n64# 0.341152f
C314 g3_inv a_161_n1258# 2.83e-19
C315 a_n13_n1158# a_34_n1189# 0.059344f
C316 p2 a_94_n825# 0.069367f
C317 b2 a2 0.626439f
C318 gnd a_247_n251# 1.36e-19
C319 in4_NAND5 in5_NAND5 0.668932f
C320 a_n13_n541# gnd 0.180335f
C321 g1 c0 0.203571f
C322 a_94_n1118# gnd 1.36e-19
C323 w_49_n36# a_133_n10# 0.248779f
C324 g1 gnd 0.182019f
C325 s1 gnd 0.103118f
C326 vdd a_82_n1024# 1.533079f
C327 a_n6_n470# b0 1.7e-19
C328 b1 a1 0.626439f
C329 a_82_n608# c2 0.106322f
C330 in1_NAND3 gnd 0.001614f
C331 in1_NAND4 out_NAND4 0.001572f
C332 a_116_n1412# gnd 0.056049f
C333 vdd g2 0.227839f
C334 c4 vdd 1.35816f
C335 g1 g1_inv 0.063031f
C336 p1 a_82_n504# 0.069367f
C337 g0_inv vdd 0.497506f
C338 in2_NAND4 in3_NAND4 0.338625f
C339 in1_NAND4 in4_NAND4 0.007681f
C340 g0 a_114_n1241# 1.7e-19
C341 vdd a_94_n825# 0.683378f
C342 a_34_n572# p1 0.060435f
C343 a_169_n498# a_216_n473# 0.059344f
C344 c0 a_82_n1024# 0.007111f
C345 in3_NAND3 a_65_n217# 2.83e-19
C346 vdd a2 0.046605f
C347 gnd a_82_n1024# 0.013419f
C348 in5_NAND5 vdd 0.020472f
C349 gnd g2 0.123737f
C350 a_100_n1287# p3 0.068884f
C351 a_197_n1258# gnd 1.36e-19
C352 c4 gnd 2.27e-20
C353 a1 vdd 0.046605f
C354 a_197_n378# s0 0.059344f
C355 c0 g0_inv 0.017409f
C356 g0_inv gnd 0.317334f
C357 a_94_n825# gnd 0.012692f
C358 a_216_n473# vdd 0.467651f
C359 in1_NAND2 in2_NAND2 0.174076f
C360 a_n13_n1158# b3 1.51355f
C361 g0_inv a0 0.036296f
C362 g3_inv p2 0.013429f
C363 a_88_n704# a_94_n825# 0.352371f
C364 a2 gnd 0.001614f
C365 in5_NAND5 gnd 0.0559f
C366 a_90_n1164# p1 0.00699f
C367 a_212_n29# in1_xor 1.51355f
C368 g1 g0 0.022143f
C369 in2_NAND2 vdd 0.020473f
C370 a_100_n1287# a_110_n1392# 1.65824f
C371 in1_xor in2_xor 0.424419f
C372 a3 g3_inv 0.036296f
C373 w_49_n36# out_ff 0.22794f
C374 in4_NAND4 out_NAND4 0.071017f
C375 in3_NAND5 in5_NAND5 0.007681f
C376 gnd a_163_n234# 1.36e-19
C377 a1 gnd 0.001614f
C378 a_161_n1258# gnd 1.36e-19
C379 a_82_n1118# gnd 1.36e-19
C380 w_49_n36# a_98_n10# 0.272577f
C381 p0 a_82_n504# 0.106322f
C382 a_148_n564# gnd 1.36e-19
C383 a_216_n473# gnd 0.262811f
C384 a_151_n725# c2 1.51355f
C385 p1 m2_67_n574# 5.76e-19
C386 a_82_n504# c2 0.036296f
C387 g1_inv a1 0.036296f
C388 in2_NAND2 gnd 0.0559f
C389 vdd s3 0.214182f
C390 g3_inv vdd 0.493348f
C391 a_82_n651# p1 1.7e-19
C392 a_148_n564# g1_inv 1.7e-19
C393 a_73_n357# vdd 0.468641f
C394 in1_NAND4 in3_NAND4 0.007278f
C395 g2_inv a_182_n845# 1.7e-19
C396 vdd a_n13_n352# 0.31023f
C397 a_268_n808# s3 0.059344f
C398 vdd b2 0.067865f
C399 in4_NAND5 vdd 0.020472f
C400 gnd a_94_n972# 1.36e-19
C401 in_ff a_51_n72# 0.056598f
C402 a_118_n1118# gnd 1.36e-19
C403 g0_inv g0 0.139333f
C404 g0 a_94_n825# 0.106322f
C405 p2 vdd 1.141294f
C406 gnd s3 0.103118f
C407 a_90_n1164# p3 0.010538f
C408 b1 vdd 0.067865f
C409 g3_inv gnd 0.810813f
C410 c0 a_73_n357# 0.163729f
C411 a3 vdd 0.046605f
C412 a_73_n357# gnd 0.001637f
C413 p2 a_106_n885# 1.7e-19
C414 c3 g2_inv 0.071017f
C415 a_112_n781# gnd 1.36e-19
C416 p3 a_112_n1347# 1.7e-19
C417 gnd a_110_n1435# 1.36e-19
C418 a_169_n498# vdd 0.31015f
C419 p0 a_150_n403# 1.51355f
C420 g0_inv b0 0.153419f
C421 a_100_n1287# g1 0.036296f
C422 a_n13_n777# a_34_n808# 0.059344f
C423 p3 c3 0.672902f
C424 b2 gnd 0.114196f
C425 gnd a_n13_n352# 0.180335f
C426 in4_NAND5 gnd 8.87e-19
C427 in1_NAND2 vdd 0.020614f
C428 p2 c0 0.226466f
C429 a_90_n1164# a_110_n1392# 0.007278f
C430 w_49_n36# a_62_n64# 0.020872f
C431 p2 gnd 0.179628f
C432 a0 a_n13_n352# 0.90085f
C433 in2_NAND5 in5_NAND5 0.007681f
C434 in3_NAND5 in4_NAND5 0.503577f
C435 gnd a_151_n234# 1.36e-19
C436 in3_NAND4 out_NAND4 0.010538f
C437 p1 g2_inv 0.001792f
C438 b1 gnd 0.114196f
C439 a3 gnd 0.001614f
C440 a_n6_n1276# gnd 1.36e-19
C441 w_49_n36# clk 0.069031f
C442 p2 a_88_n704# 0.001572f
C443 p0 p1 1.37465f
C444 a_136_n564# gnd 1.36e-19
C445 p1 p3 0.594173f
C446 in3_NAND4 in4_NAND4 0.50398f
C447 a_169_n498# gnd 0.180335f
C448 p2 g1_inv 0.701046f
C449 g1_inv b1 0.153419f
C450 in1_NAND2 gnd 0.001614f
C451 in2_NAND2 a_n6_n200# 1.7e-19
C452 in3_NAND3 out_NAND3 0.069367f
C453 vdd a_268_n808# 0.467651f
C454 a_100_n1287# a_82_n1024# 0.007278f
C455 a_34_n572# a_n13_n541# 0.059344f
C456 a_136_n564# g1_inv 2.83e-19
C457 c0 vdd 0.203741f
C458 vdd gnd 0.85308f
C459 g3_inv a_173_n1258# 2.83e-19
C460 a_100_n1287# c4 0.007111f
C461 g3_inv g0 8.39e-22
C462 g2_inv a_170_n845# 2.83e-19
C463 vdd a_88_n704# 1.041384f
C464 gnd a_106_n885# 1.36e-19
C465 in3_NAND5 vdd 0.020472f
C466 vdd a0 0.046605f
C467 g0_inv a_108_n400# 1.7e-19
C468 s2 vdd 0.214182f
C469 gnd a_268_n808# 0.262811f
C470 a_34_n1189# p3 0.059344f
C471 g1_inv vdd 0.489081f
C472 in2_NAND3 in3_NAND3 0.339028f
C473 p0 g2_inv 0.009794f
C474 c0 gnd 0.915614f
C475 p2 a_94_n885# 2.83e-19
C476 p3 g2_inv 0.003344f
C477 c3 a_94_n929# 0.010538f
C478 a_100_n781# gnd 1.36e-19
C479 a_133_n50# a_51_n72# 1.36e-19
C480 p2 g0 0.60512f
C481 c0 a_88_n704# 0.00699f
C482 a_34_n383# a_n13_n352# 0.059344f
C483 p0 p3 0.006063f
C484 gnd a0 0.001614f
C485 a_88_n704# gnd 0.001637f
C486 in5_NAND5 out_NAND5 0.071424f
C487 in3_NAND5 gnd 8.87e-19
C488 out_xor vdd 0.214182f
C489 m2_67_n574# 0 0.08181f
C490 m2_37_n508# 0 0.082199f
C491 gnd 0 5.822654f **FLOATING
C492 a_116_n1412# 0 0.875719f **FLOATING
C493 g3 0 0.067079f **FLOATING
C494 c4 0 0.364336f **FLOATING
C495 g3_inv 0 1.44395f **FLOATING
C496 a_110_n1392# 0 1.05172f **FLOATING
C497 a_100_n1287# 0 0.747773f **FLOATING
C498 a_90_n1164# 0 0.600617f **FLOATING
C499 a_34_n1189# 0 0.225278f **FLOATING
C500 a_n13_n1158# 0 0.429392f **FLOATING
C501 a3 0 0.632398f **FLOATING
C502 b3 0 1.39887f **FLOATING
C503 a_82_n1024# 0 0.84293f **FLOATING
C504 g2 0 0.078517f **FLOATING
C505 s3 0 0.098366f **FLOATING
C506 a_268_n808# 0 0.225278f **FLOATING
C507 a_221_n777# 0 0.429392f **FLOATING
C508 g2_inv 0 1.66541f **FLOATING
C509 a_94_n929# 0 0.74302f **FLOATING
C510 a_94_n825# 0 0.72596f **FLOATING
C511 a_34_n808# 0 0.225278f **FLOATING
C512 c3 0 0.47077f **FLOATING
C513 p3 0 3.16721f **FLOATING
C514 a_n13_n777# 0 0.429392f **FLOATING
C515 a2 0 0.632398f **FLOATING
C516 b2 0 1.39887f **FLOATING
C517 a_88_n704# 0 0.610966f **FLOATING
C518 p2 0 3.54345f **FLOATING
C519 s2 0 0.098366f **FLOATING
C520 a_198_n700# 0 0.225278f **FLOATING
C521 a_151_n725# 0 0.400729f **FLOATING
C522 g1 0 7.93276f **FLOATING
C523 a_34_n572# 0 0.225278f **FLOATING
C524 c2 0 0.845223f **FLOATING
C525 a_n13_n541# 0 0.429392f **FLOATING
C526 a1 0 0.632398f **FLOATING
C527 b1 0 1.39887f **FLOATING
C528 g1_inv 0 1.16183f **FLOATING
C529 a_82_n608# 0 0.614698f **FLOATING
C530 a_82_n504# 0 0.496897f **FLOATING
C531 p1 0 5.02911f **FLOATING
C532 s1 0 0.098366f **FLOATING
C533 a_216_n473# 0 0.225278f **FLOATING
C534 a_169_n498# 0 0.405811f **FLOATING
C535 g0 0 3.77874f **FLOATING
C536 s0 0 0.098366f **FLOATING
C537 c1 0 0.767831f **FLOATING
C538 g0_inv 0 2.34788f **FLOATING
C539 a_73_n357# 0 0.356625f **FLOATING
C540 c0 0 7.29956f **FLOATING
C541 a_34_n383# 0 0.225278f **FLOATING
C542 a_197_n378# 0 0.225278f **FLOATING
C543 a_150_n403# 0 0.373172f **FLOATING
C544 p0 0 2.57423f **FLOATING
C545 a_n13_n352# 0 0.429392f **FLOATING
C546 a0 0 0.632398f **FLOATING
C547 b0 0 1.39887f **FLOATING
C548 out_NAND5 0 0.364336f **FLOATING
C549 out_NAND4 0 0.293488f **FLOATING
C550 out_NAND3 0 0.275637f **FLOATING
C551 out_NAND2 0 0.154398f **FLOATING
C552 in5_NAND5 0 0.452425f **FLOATING
C553 in4_NAND5 0 0.38217f **FLOATING
C554 in3_NAND5 0 0.369292f **FLOATING
C555 in2_NAND5 0 0.356414f **FLOATING
C556 in1_NAND5 0 0.346357f **FLOATING
C557 in4_NAND4 0 0.38724f **FLOATING
C558 in3_NAND4 0 0.328622f **FLOATING
C559 in2_NAND4 0 0.315744f **FLOATING
C560 in1_NAND4 0 0.305687f **FLOATING
C561 in3_NAND3 0 0.322054f **FLOATING
C562 in2_NAND3 0 0.268145f **FLOATING
C563 in1_NAND3 0 0.26109f **FLOATING
C564 in2_NAND2 0 0.24994f **FLOATING
C565 in1_NAND2 0 0.22042f **FLOATING
C566 out_xor 0 0.098366f **FLOATING
C567 a_259_n60# 0 0.225278f **FLOATING
C568 a_212_n29# 0 0.429392f **FLOATING
C569 a_51_n72# 0 0.542627f **FLOATING
C570 out_ff 0 0.094438f **FLOATING
C571 a_62_n64# 0 0.323967f **FLOATING
C572 out_inv 0 0.098366f **FLOATING
C573 in_inv 0 0.194444f **FLOATING
C574 in2_xor 0 0.170441f **FLOATING
C575 in1_xor 0 0.266338f **FLOATING
C576 a_133_n10# 0 0.299294f **FLOATING
C577 a_98_n10# 0 0.33934f **FLOATING
C578 clk 0 1.56137f **FLOATING
C579 in_ff 0 0.222447f **FLOATING
C580 vdd 0 83.2702f **FLOATING
C581 w_49_n36# 0 5.96533f **FLOATING
