magic
tech scmos
timestamp 1732015174
<< nwell >>
rect -26 -25 -2 14
rect 49 -16 172 23
rect 206 -1 246 24
rect 49 -36 85 -16
rect 206 -35 286 -1
rect 246 -40 286 -35
rect -19 -163 17 -124
rect 52 -163 100 -124
rect 126 -163 186 -124
rect 234 -163 306 -124
rect -19 -324 21 -299
rect -19 -358 131 -324
rect 184 -357 224 -352
rect 21 -363 131 -358
rect 144 -391 224 -357
rect -19 -433 33 -394
rect 144 -416 184 -391
rect 203 -452 243 -447
rect 163 -471 243 -452
rect -19 -513 21 -488
rect 69 -510 117 -471
rect 123 -486 243 -471
rect 123 -510 203 -486
rect 163 -511 203 -510
rect -19 -547 61 -513
rect 21 -552 61 -547
rect -19 -622 33 -583
rect 69 -614 105 -575
rect 75 -710 135 -671
rect 185 -679 225 -674
rect 145 -715 225 -679
rect -19 -749 21 -724
rect 145 -735 185 -715
rect -19 -783 61 -749
rect 145 -774 205 -735
rect 215 -749 255 -724
rect 215 -783 295 -749
rect 21 -788 61 -783
rect 255 -788 295 -783
rect -19 -858 33 -819
rect 81 -831 129 -792
rect 81 -935 117 -896
rect 69 -1030 141 -991
rect -19 -1130 21 -1105
rect -19 -1164 61 -1130
rect 21 -1169 61 -1164
rect 77 -1170 137 -1131
rect 148 -1170 220 -1131
rect -19 -1239 33 -1200
rect 87 -1293 135 -1253
rect 97 -1398 133 -1359
<< ntransistor >>
rect -15 -45 -13 -35
rect 96 -50 98 -30
rect 108 -50 110 -30
rect 131 -50 133 -30
rect 143 -50 145 -30
rect 159 -36 161 -26
rect 60 -64 62 -54
rect 217 -60 219 -50
rect 257 -60 259 -50
rect 273 -60 275 -50
rect -8 -200 -6 -180
rect 4 -200 6 -180
rect 63 -217 65 -187
rect 75 -217 77 -187
rect 87 -217 89 -187
rect 137 -234 139 -194
rect 149 -234 151 -194
rect 161 -234 163 -194
rect 173 -234 175 -194
rect 245 -251 247 -201
rect 257 -251 259 -201
rect 269 -251 271 -201
rect 281 -251 283 -201
rect 293 -251 295 -201
rect 155 -342 157 -332
rect 195 -342 197 -332
rect 211 -342 213 -332
rect -8 -383 -6 -373
rect 32 -383 34 -373
rect 48 -383 50 -373
rect 71 -400 73 -380
rect 83 -400 85 -380
rect 106 -400 108 -380
rect 118 -400 120 -380
rect 174 -437 176 -427
rect 214 -437 216 -427
rect 230 -437 232 -427
rect -8 -470 -6 -450
rect 4 -470 6 -450
rect 20 -453 22 -443
rect -8 -572 -6 -562
rect 32 -572 34 -562
rect 48 -572 50 -562
rect 80 -564 82 -534
rect 92 -564 94 -534
rect 104 -564 106 -534
rect 134 -564 136 -534
rect 146 -564 148 -534
rect 158 -564 160 -534
rect -8 -659 -6 -639
rect 4 -659 6 -639
rect 20 -642 22 -632
rect 80 -651 82 -631
rect 92 -651 94 -631
rect 156 -664 158 -654
rect 196 -664 198 -654
rect 212 -664 214 -654
rect 86 -781 88 -741
rect 98 -781 100 -741
rect 110 -781 112 -741
rect 122 -781 124 -741
rect -8 -808 -6 -798
rect 32 -808 34 -798
rect 48 -808 50 -798
rect 156 -845 158 -805
rect 168 -845 170 -805
rect 180 -845 182 -805
rect 192 -845 194 -805
rect 226 -808 228 -798
rect 266 -808 268 -798
rect 282 -808 284 -798
rect -8 -895 -6 -875
rect 4 -895 6 -875
rect 20 -878 22 -868
rect 92 -885 94 -855
rect 104 -885 106 -855
rect 116 -885 118 -855
rect 92 -972 94 -952
rect 104 -972 106 -952
rect 80 -1118 82 -1068
rect 92 -1118 94 -1068
rect 104 -1118 106 -1068
rect 116 -1118 118 -1068
rect 128 -1118 130 -1068
rect -8 -1189 -6 -1179
rect 32 -1189 34 -1179
rect 48 -1189 50 -1179
rect 88 -1241 90 -1201
rect 100 -1241 102 -1201
rect 112 -1241 114 -1201
rect 124 -1241 126 -1201
rect -8 -1276 -6 -1256
rect 4 -1276 6 -1256
rect 20 -1259 22 -1249
rect 159 -1258 161 -1208
rect 171 -1258 173 -1208
rect 183 -1258 185 -1208
rect 195 -1258 197 -1208
rect 207 -1258 209 -1208
rect 98 -1347 100 -1317
rect 110 -1347 112 -1317
rect 122 -1347 124 -1317
rect 108 -1435 110 -1415
rect 120 -1435 122 -1415
<< ptransistor >>
rect -15 -19 -13 1
rect 60 -30 62 10
rect 72 -30 74 10
rect 96 -10 98 10
rect 131 -10 133 10
rect 159 -10 161 10
rect 217 -29 219 11
rect 233 -29 235 11
rect 257 -34 259 -14
rect 273 -34 275 -14
rect -8 -157 -6 -137
rect 4 -157 6 -137
rect 63 -157 65 -137
rect 75 -157 77 -137
rect 87 -157 89 -137
rect 137 -157 139 -137
rect 149 -157 151 -137
rect 161 -157 163 -137
rect 173 -157 175 -137
rect 245 -157 247 -137
rect 257 -157 259 -137
rect 269 -157 271 -137
rect 281 -157 283 -137
rect 293 -157 295 -137
rect -8 -352 -6 -312
rect 8 -352 10 -312
rect 32 -357 34 -337
rect 48 -357 50 -337
rect 71 -357 73 -337
rect 83 -357 85 -337
rect 106 -357 108 -337
rect 118 -357 120 -337
rect 155 -403 157 -363
rect 171 -403 173 -363
rect 195 -378 197 -358
rect 211 -378 213 -358
rect -8 -427 -6 -407
rect 4 -427 6 -407
rect 20 -427 22 -407
rect -8 -541 -6 -501
rect 8 -541 10 -501
rect 80 -504 82 -484
rect 92 -504 94 -484
rect 104 -504 106 -484
rect 134 -504 136 -484
rect 146 -504 148 -484
rect 158 -504 160 -484
rect 174 -498 176 -458
rect 190 -498 192 -458
rect 214 -473 216 -453
rect 230 -473 232 -453
rect 32 -546 34 -526
rect 48 -546 50 -526
rect -8 -616 -6 -596
rect 4 -616 6 -596
rect 20 -616 22 -596
rect 80 -608 82 -588
rect 92 -608 94 -588
rect 86 -704 88 -684
rect 98 -704 100 -684
rect 110 -704 112 -684
rect 122 -704 124 -684
rect -8 -777 -6 -737
rect 8 -777 10 -737
rect 156 -725 158 -685
rect 172 -725 174 -685
rect 196 -700 198 -680
rect 212 -700 214 -680
rect 32 -782 34 -762
rect 48 -782 50 -762
rect 156 -768 158 -748
rect 168 -768 170 -748
rect 180 -768 182 -748
rect 192 -768 194 -748
rect 226 -777 228 -737
rect 242 -777 244 -737
rect 266 -782 268 -762
rect 282 -782 284 -762
rect 92 -825 94 -805
rect 104 -825 106 -805
rect 116 -825 118 -805
rect -8 -852 -6 -832
rect 4 -852 6 -832
rect 20 -852 22 -832
rect 92 -929 94 -909
rect 104 -929 106 -909
rect 80 -1024 82 -1004
rect 92 -1024 94 -1004
rect 104 -1024 106 -1004
rect 116 -1024 118 -1004
rect 128 -1024 130 -1004
rect -8 -1158 -6 -1118
rect 8 -1158 10 -1118
rect 32 -1163 34 -1143
rect 48 -1163 50 -1143
rect 88 -1164 90 -1144
rect 100 -1164 102 -1144
rect 112 -1164 114 -1144
rect 124 -1164 126 -1144
rect 159 -1164 161 -1144
rect 171 -1164 173 -1144
rect 183 -1164 185 -1144
rect 195 -1164 197 -1144
rect 207 -1164 209 -1144
rect -8 -1233 -6 -1213
rect 4 -1233 6 -1213
rect 20 -1233 22 -1213
rect 98 -1287 100 -1267
rect 110 -1287 112 -1267
rect 122 -1287 124 -1267
rect 108 -1392 110 -1372
rect 120 -1392 122 -1372
<< ndiffusion >>
rect -16 -45 -15 -35
rect -13 -45 -12 -35
rect 95 -50 96 -30
rect 98 -50 108 -30
rect 110 -50 111 -30
rect 130 -50 131 -30
rect 133 -50 143 -30
rect 145 -50 146 -30
rect 158 -36 159 -26
rect 161 -36 162 -26
rect 59 -64 60 -54
rect 62 -64 63 -54
rect 216 -60 217 -50
rect 219 -60 220 -50
rect 256 -60 257 -50
rect 259 -60 260 -50
rect 272 -60 273 -50
rect 275 -60 276 -50
rect -9 -200 -8 -180
rect -6 -200 4 -180
rect 6 -200 7 -180
rect 62 -217 63 -187
rect 65 -217 75 -187
rect 77 -217 87 -187
rect 89 -217 90 -187
rect 136 -234 137 -194
rect 139 -234 149 -194
rect 151 -234 161 -194
rect 163 -234 173 -194
rect 175 -234 176 -194
rect 244 -251 245 -201
rect 247 -251 257 -201
rect 259 -251 269 -201
rect 271 -251 281 -201
rect 283 -251 293 -201
rect 295 -251 296 -201
rect 154 -342 155 -332
rect 157 -342 158 -332
rect 194 -342 195 -332
rect 197 -342 198 -332
rect 210 -342 211 -332
rect 213 -342 214 -332
rect -9 -383 -8 -373
rect -6 -383 -5 -373
rect 31 -383 32 -373
rect 34 -383 35 -373
rect 47 -383 48 -373
rect 50 -383 51 -373
rect 70 -400 71 -380
rect 73 -400 83 -380
rect 85 -400 86 -380
rect 105 -400 106 -380
rect 108 -400 118 -380
rect 120 -400 121 -380
rect 173 -437 174 -427
rect 176 -437 177 -427
rect 213 -437 214 -427
rect 216 -437 217 -427
rect 229 -437 230 -427
rect 232 -437 233 -427
rect -9 -470 -8 -450
rect -6 -470 4 -450
rect 6 -470 7 -450
rect 19 -453 20 -443
rect 22 -453 23 -443
rect -9 -572 -8 -562
rect -6 -572 -5 -562
rect 31 -572 32 -562
rect 34 -572 35 -562
rect 47 -572 48 -562
rect 50 -572 51 -562
rect 79 -564 80 -534
rect 82 -564 92 -534
rect 94 -564 104 -534
rect 106 -564 107 -534
rect 133 -564 134 -534
rect 136 -564 146 -534
rect 148 -564 158 -534
rect 160 -564 161 -534
rect -9 -659 -8 -639
rect -6 -659 4 -639
rect 6 -659 7 -639
rect 19 -642 20 -632
rect 22 -642 23 -632
rect 79 -651 80 -631
rect 82 -651 92 -631
rect 94 -651 95 -631
rect 155 -664 156 -654
rect 158 -664 159 -654
rect 195 -664 196 -654
rect 198 -664 199 -654
rect 211 -664 212 -654
rect 214 -664 215 -654
rect 85 -781 86 -741
rect 88 -781 98 -741
rect 100 -781 110 -741
rect 112 -781 122 -741
rect 124 -781 125 -741
rect -9 -808 -8 -798
rect -6 -808 -5 -798
rect 31 -808 32 -798
rect 34 -808 35 -798
rect 47 -808 48 -798
rect 50 -808 51 -798
rect 155 -845 156 -805
rect 158 -845 168 -805
rect 170 -845 180 -805
rect 182 -845 192 -805
rect 194 -845 195 -805
rect 225 -808 226 -798
rect 228 -808 229 -798
rect 265 -808 266 -798
rect 268 -808 269 -798
rect 281 -808 282 -798
rect 284 -808 285 -798
rect -9 -895 -8 -875
rect -6 -895 4 -875
rect 6 -895 7 -875
rect 19 -878 20 -868
rect 22 -878 23 -868
rect 91 -885 92 -855
rect 94 -885 104 -855
rect 106 -885 116 -855
rect 118 -885 119 -855
rect 91 -972 92 -952
rect 94 -972 104 -952
rect 106 -972 107 -952
rect 79 -1118 80 -1068
rect 82 -1118 92 -1068
rect 94 -1118 104 -1068
rect 106 -1118 116 -1068
rect 118 -1118 128 -1068
rect 130 -1118 131 -1068
rect -9 -1189 -8 -1179
rect -6 -1189 -5 -1179
rect 31 -1189 32 -1179
rect 34 -1189 35 -1179
rect 47 -1189 48 -1179
rect 50 -1189 51 -1179
rect 87 -1241 88 -1201
rect 90 -1241 100 -1201
rect 102 -1241 112 -1201
rect 114 -1241 124 -1201
rect 126 -1241 127 -1201
rect -9 -1276 -8 -1256
rect -6 -1276 4 -1256
rect 6 -1276 7 -1256
rect 19 -1259 20 -1249
rect 22 -1259 23 -1249
rect 158 -1258 159 -1208
rect 161 -1258 171 -1208
rect 173 -1258 183 -1208
rect 185 -1258 195 -1208
rect 197 -1258 207 -1208
rect 209 -1258 210 -1208
rect 97 -1347 98 -1317
rect 100 -1347 110 -1317
rect 112 -1347 122 -1317
rect 124 -1347 125 -1317
rect 107 -1435 108 -1415
rect 110 -1435 120 -1415
rect 122 -1435 123 -1415
<< pdiffusion >>
rect -16 -19 -15 1
rect -13 -19 -12 1
rect 59 -30 60 10
rect 62 -30 72 10
rect 74 -30 75 10
rect 95 -10 96 10
rect 98 -10 99 10
rect 130 -10 131 10
rect 133 -10 134 10
rect 158 -10 159 10
rect 161 -10 162 10
rect 216 -29 217 11
rect 219 -29 220 11
rect 232 -29 233 11
rect 235 -29 236 11
rect 256 -34 257 -14
rect 259 -34 260 -14
rect 272 -34 273 -14
rect 275 -34 276 -14
rect -9 -157 -8 -137
rect -6 -157 -5 -137
rect 3 -157 4 -137
rect 6 -157 7 -137
rect 62 -157 63 -137
rect 65 -157 66 -137
rect 74 -157 75 -137
rect 77 -157 78 -137
rect 86 -157 87 -137
rect 89 -157 90 -137
rect 136 -157 137 -137
rect 139 -157 140 -137
rect 148 -157 149 -137
rect 151 -157 152 -137
rect 160 -157 161 -137
rect 163 -157 164 -137
rect 172 -157 173 -137
rect 175 -157 176 -137
rect 244 -157 245 -137
rect 247 -157 248 -137
rect 256 -157 257 -137
rect 259 -157 260 -137
rect 268 -157 269 -137
rect 271 -157 272 -137
rect 280 -157 281 -137
rect 283 -157 284 -137
rect 292 -157 293 -137
rect 295 -157 296 -137
rect -9 -352 -8 -312
rect -6 -352 -5 -312
rect 7 -352 8 -312
rect 10 -352 11 -312
rect 31 -357 32 -337
rect 34 -357 35 -337
rect 47 -357 48 -337
rect 50 -357 51 -337
rect 70 -357 71 -337
rect 73 -357 74 -337
rect 82 -357 83 -337
rect 85 -357 86 -337
rect 105 -357 106 -337
rect 108 -357 109 -337
rect 117 -357 118 -337
rect 120 -357 121 -337
rect 154 -403 155 -363
rect 157 -403 158 -363
rect 170 -403 171 -363
rect 173 -403 174 -363
rect 194 -378 195 -358
rect 197 -378 198 -358
rect 210 -378 211 -358
rect 213 -378 214 -358
rect -9 -427 -8 -407
rect -6 -427 -5 -407
rect 3 -427 4 -407
rect 6 -427 7 -407
rect 19 -427 20 -407
rect 22 -427 23 -407
rect -9 -541 -8 -501
rect -6 -541 -5 -501
rect 7 -541 8 -501
rect 10 -541 11 -501
rect 79 -504 80 -484
rect 82 -504 83 -484
rect 91 -504 92 -484
rect 94 -504 95 -484
rect 103 -504 104 -484
rect 106 -504 107 -484
rect 133 -504 134 -484
rect 136 -504 137 -484
rect 145 -504 146 -484
rect 148 -504 149 -484
rect 157 -504 158 -484
rect 160 -504 161 -484
rect 173 -498 174 -458
rect 176 -498 177 -458
rect 189 -498 190 -458
rect 192 -498 193 -458
rect 213 -473 214 -453
rect 216 -473 217 -453
rect 229 -473 230 -453
rect 232 -473 233 -453
rect 31 -546 32 -526
rect 34 -546 35 -526
rect 47 -546 48 -526
rect 50 -546 51 -526
rect -9 -616 -8 -596
rect -6 -616 -5 -596
rect 3 -616 4 -596
rect 6 -616 7 -596
rect 19 -616 20 -596
rect 22 -616 23 -596
rect 79 -608 80 -588
rect 82 -608 83 -588
rect 91 -608 92 -588
rect 94 -608 95 -588
rect 85 -704 86 -684
rect 88 -704 89 -684
rect 97 -704 98 -684
rect 100 -704 101 -684
rect 109 -704 110 -684
rect 112 -704 113 -684
rect 121 -704 122 -684
rect 124 -704 125 -684
rect -9 -777 -8 -737
rect -6 -777 -5 -737
rect 7 -777 8 -737
rect 10 -777 11 -737
rect 155 -725 156 -685
rect 158 -725 159 -685
rect 171 -725 172 -685
rect 174 -725 175 -685
rect 195 -700 196 -680
rect 198 -700 199 -680
rect 211 -700 212 -680
rect 214 -700 215 -680
rect 31 -782 32 -762
rect 34 -782 35 -762
rect 47 -782 48 -762
rect 50 -782 51 -762
rect 155 -768 156 -748
rect 158 -768 159 -748
rect 167 -768 168 -748
rect 170 -768 171 -748
rect 179 -768 180 -748
rect 182 -768 183 -748
rect 191 -768 192 -748
rect 194 -768 195 -748
rect 225 -777 226 -737
rect 228 -777 229 -737
rect 241 -777 242 -737
rect 244 -777 245 -737
rect 265 -782 266 -762
rect 268 -782 269 -762
rect 281 -782 282 -762
rect 284 -782 285 -762
rect 91 -825 92 -805
rect 94 -825 95 -805
rect 103 -825 104 -805
rect 106 -825 107 -805
rect 115 -825 116 -805
rect 118 -825 119 -805
rect -9 -852 -8 -832
rect -6 -852 -5 -832
rect 3 -852 4 -832
rect 6 -852 7 -832
rect 19 -852 20 -832
rect 22 -852 23 -832
rect 91 -929 92 -909
rect 94 -929 95 -909
rect 103 -929 104 -909
rect 106 -929 107 -909
rect 79 -1024 80 -1004
rect 82 -1024 83 -1004
rect 91 -1024 92 -1004
rect 94 -1024 95 -1004
rect 103 -1024 104 -1004
rect 106 -1024 107 -1004
rect 115 -1024 116 -1004
rect 118 -1024 119 -1004
rect 127 -1024 128 -1004
rect 130 -1024 131 -1004
rect -9 -1158 -8 -1118
rect -6 -1158 -5 -1118
rect 7 -1158 8 -1118
rect 10 -1158 11 -1118
rect 31 -1163 32 -1143
rect 34 -1163 35 -1143
rect 47 -1163 48 -1143
rect 50 -1163 51 -1143
rect 87 -1164 88 -1144
rect 90 -1164 91 -1144
rect 99 -1164 100 -1144
rect 102 -1164 103 -1144
rect 111 -1164 112 -1144
rect 114 -1164 115 -1144
rect 123 -1164 124 -1144
rect 126 -1164 127 -1144
rect 158 -1164 159 -1144
rect 161 -1164 162 -1144
rect 170 -1164 171 -1144
rect 173 -1164 174 -1144
rect 182 -1164 183 -1144
rect 185 -1164 186 -1144
rect 194 -1164 195 -1144
rect 197 -1164 198 -1144
rect 206 -1164 207 -1144
rect 209 -1164 210 -1144
rect -9 -1233 -8 -1213
rect -6 -1233 -5 -1213
rect 3 -1233 4 -1213
rect 6 -1233 7 -1213
rect 19 -1233 20 -1213
rect 22 -1233 23 -1213
rect 97 -1287 98 -1267
rect 100 -1287 101 -1267
rect 109 -1287 110 -1267
rect 112 -1287 113 -1267
rect 121 -1287 122 -1267
rect 124 -1287 125 -1267
rect 107 -1392 108 -1372
rect 110 -1392 111 -1372
rect 119 -1392 120 -1372
rect 122 -1392 123 -1372
<< ndcontact >>
rect -20 -45 -16 -35
rect -12 -45 -8 -35
rect 91 -50 95 -30
rect 111 -50 115 -30
rect 126 -50 130 -30
rect 146 -50 150 -30
rect 154 -36 158 -26
rect 162 -36 166 -26
rect 55 -64 59 -54
rect 63 -64 67 -54
rect 212 -60 216 -50
rect 220 -60 224 -50
rect 252 -60 256 -50
rect 260 -60 264 -50
rect 268 -60 272 -50
rect 276 -60 280 -50
rect -13 -200 -9 -180
rect 7 -200 11 -180
rect 58 -217 62 -187
rect 90 -217 94 -187
rect 132 -234 136 -194
rect 176 -234 180 -194
rect 240 -251 244 -201
rect 296 -251 300 -201
rect 150 -342 154 -332
rect 158 -342 162 -332
rect 190 -342 194 -332
rect 198 -342 202 -332
rect 206 -342 210 -332
rect 214 -342 218 -332
rect -13 -383 -9 -373
rect -5 -383 -1 -373
rect 27 -383 31 -373
rect 35 -383 39 -373
rect 43 -383 47 -373
rect 51 -383 55 -373
rect 66 -400 70 -380
rect 86 -400 90 -380
rect 101 -400 105 -380
rect 121 -400 125 -380
rect 169 -437 173 -427
rect 177 -437 181 -427
rect 209 -437 213 -427
rect 217 -437 221 -427
rect 225 -437 229 -427
rect 233 -437 237 -427
rect -13 -470 -9 -450
rect 7 -470 11 -450
rect 15 -453 19 -443
rect 23 -453 27 -443
rect -13 -572 -9 -562
rect -5 -572 -1 -562
rect 27 -572 31 -562
rect 35 -572 39 -562
rect 43 -572 47 -562
rect 51 -572 55 -562
rect 75 -564 79 -534
rect 107 -564 111 -534
rect 129 -564 133 -534
rect 161 -564 165 -534
rect -13 -659 -9 -639
rect 7 -659 11 -639
rect 15 -642 19 -632
rect 23 -642 27 -632
rect 75 -651 79 -631
rect 95 -651 99 -631
rect 151 -664 155 -654
rect 159 -664 163 -654
rect 191 -664 195 -654
rect 199 -664 203 -654
rect 207 -664 211 -654
rect 215 -664 219 -654
rect 81 -781 85 -741
rect 125 -781 129 -741
rect -13 -808 -9 -798
rect -5 -808 -1 -798
rect 27 -808 31 -798
rect 35 -808 39 -798
rect 43 -808 47 -798
rect 51 -808 55 -798
rect 151 -845 155 -805
rect 195 -845 199 -805
rect 221 -808 225 -798
rect 229 -808 233 -798
rect 261 -808 265 -798
rect 269 -808 273 -798
rect 277 -808 281 -798
rect 285 -808 289 -798
rect -13 -895 -9 -875
rect 7 -895 11 -875
rect 15 -878 19 -868
rect 23 -878 27 -868
rect 87 -885 91 -855
rect 119 -885 123 -855
rect 87 -972 91 -952
rect 107 -972 111 -952
rect 75 -1118 79 -1068
rect 131 -1118 135 -1068
rect -13 -1189 -9 -1179
rect -5 -1189 -1 -1179
rect 27 -1189 31 -1179
rect 35 -1189 39 -1179
rect 43 -1189 47 -1179
rect 51 -1189 55 -1179
rect 83 -1241 87 -1201
rect 127 -1241 131 -1201
rect -13 -1276 -9 -1256
rect 7 -1276 11 -1256
rect 15 -1259 19 -1249
rect 23 -1259 27 -1249
rect 154 -1258 158 -1208
rect 210 -1258 214 -1208
rect 93 -1347 97 -1317
rect 125 -1347 129 -1317
rect 103 -1435 107 -1415
rect 123 -1435 127 -1415
<< pdcontact >>
rect -20 -19 -16 1
rect -12 -19 -8 1
rect 55 -30 59 10
rect 75 -30 79 10
rect 91 -10 95 10
rect 99 -10 103 10
rect 126 -10 130 10
rect 134 -10 138 10
rect 154 -10 158 10
rect 162 -10 166 10
rect 212 -29 216 11
rect 220 -29 224 11
rect 228 -29 232 11
rect 236 -29 240 11
rect 252 -34 256 -14
rect 260 -34 264 -14
rect 268 -34 272 -14
rect 276 -34 280 -14
rect -13 -157 -9 -137
rect -5 -157 3 -137
rect 7 -157 11 -137
rect 58 -157 62 -137
rect 66 -157 74 -137
rect 78 -157 86 -137
rect 90 -157 94 -137
rect 132 -157 136 -137
rect 140 -157 148 -137
rect 152 -157 160 -137
rect 164 -157 172 -137
rect 176 -157 180 -137
rect 240 -157 244 -137
rect 248 -157 256 -137
rect 260 -157 268 -137
rect 272 -157 280 -137
rect 284 -157 292 -137
rect 296 -157 300 -137
rect -13 -352 -9 -312
rect -5 -352 -1 -312
rect 3 -352 7 -312
rect 11 -352 15 -312
rect 27 -357 31 -337
rect 35 -357 39 -337
rect 43 -357 47 -337
rect 51 -357 55 -337
rect 66 -357 70 -337
rect 74 -357 82 -337
rect 86 -357 90 -337
rect 101 -357 105 -337
rect 109 -357 117 -337
rect 121 -357 125 -337
rect 150 -403 154 -363
rect 158 -403 162 -363
rect 166 -403 170 -363
rect 174 -403 178 -363
rect 190 -378 194 -358
rect 198 -378 202 -358
rect 206 -378 210 -358
rect 214 -378 218 -358
rect -13 -427 -9 -407
rect -5 -427 3 -407
rect 7 -427 11 -407
rect 15 -427 19 -407
rect 23 -427 27 -407
rect -13 -541 -9 -501
rect -5 -541 -1 -501
rect 3 -541 7 -501
rect 11 -541 15 -501
rect 75 -504 79 -484
rect 83 -504 91 -484
rect 95 -504 103 -484
rect 107 -504 111 -484
rect 129 -504 133 -484
rect 137 -504 145 -484
rect 149 -504 157 -484
rect 161 -504 165 -484
rect 169 -498 173 -458
rect 177 -498 181 -458
rect 185 -498 189 -458
rect 193 -498 197 -458
rect 209 -473 213 -453
rect 217 -473 221 -453
rect 225 -473 229 -453
rect 233 -473 237 -453
rect 27 -546 31 -526
rect 35 -546 39 -526
rect 43 -546 47 -526
rect 51 -546 55 -526
rect -13 -616 -9 -596
rect -5 -616 3 -596
rect 7 -616 11 -596
rect 15 -616 19 -596
rect 23 -616 27 -596
rect 75 -608 79 -588
rect 83 -608 91 -588
rect 95 -608 99 -588
rect 81 -704 85 -684
rect 89 -704 97 -684
rect 101 -704 109 -684
rect 113 -704 121 -684
rect 125 -704 129 -684
rect -13 -777 -9 -737
rect -5 -777 -1 -737
rect 3 -777 7 -737
rect 11 -777 15 -737
rect 151 -725 155 -685
rect 159 -725 163 -685
rect 167 -725 171 -685
rect 175 -725 179 -685
rect 191 -700 195 -680
rect 199 -700 203 -680
rect 207 -700 211 -680
rect 215 -700 219 -680
rect 27 -782 31 -762
rect 35 -782 39 -762
rect 43 -782 47 -762
rect 51 -782 55 -762
rect 151 -768 155 -748
rect 159 -768 167 -748
rect 171 -768 179 -748
rect 183 -768 191 -748
rect 195 -768 199 -748
rect 221 -777 225 -737
rect 229 -777 233 -737
rect 237 -777 241 -737
rect 245 -777 249 -737
rect 261 -782 265 -762
rect 269 -782 273 -762
rect 277 -782 281 -762
rect 285 -782 289 -762
rect 87 -825 91 -805
rect 95 -825 103 -805
rect 107 -825 115 -805
rect 119 -825 123 -805
rect -13 -852 -9 -832
rect -5 -852 3 -832
rect 7 -852 11 -832
rect 15 -852 19 -832
rect 23 -852 27 -832
rect 87 -929 91 -909
rect 95 -929 103 -909
rect 107 -929 111 -909
rect 75 -1024 79 -1004
rect 83 -1024 91 -1004
rect 95 -1024 103 -1004
rect 107 -1024 115 -1004
rect 119 -1024 127 -1004
rect 131 -1024 135 -1004
rect -13 -1158 -9 -1118
rect -5 -1158 -1 -1118
rect 3 -1158 7 -1118
rect 11 -1158 15 -1118
rect 27 -1163 31 -1143
rect 35 -1163 39 -1143
rect 43 -1163 47 -1143
rect 51 -1163 55 -1143
rect 83 -1164 87 -1144
rect 91 -1164 99 -1144
rect 103 -1164 111 -1144
rect 115 -1164 123 -1144
rect 127 -1164 131 -1144
rect 154 -1164 158 -1144
rect 162 -1164 170 -1144
rect 174 -1164 182 -1144
rect 186 -1164 194 -1144
rect 198 -1164 206 -1144
rect 210 -1164 214 -1144
rect -13 -1233 -9 -1213
rect -5 -1233 3 -1213
rect 7 -1233 11 -1213
rect 15 -1233 19 -1213
rect 23 -1233 27 -1213
rect 93 -1287 97 -1267
rect 101 -1287 109 -1267
rect 113 -1287 121 -1267
rect 125 -1287 129 -1267
rect 103 -1392 107 -1372
rect 111 -1392 119 -1372
rect 123 -1392 127 -1372
<< psubstratepcontact >>
rect -20 -53 -16 -49
rect -12 -53 -8 -49
rect 154 -44 158 -40
rect 164 -44 168 -40
rect 72 -58 76 -54
rect 87 -58 91 -54
rect 103 -58 107 -54
rect 122 -58 126 -54
rect 138 -58 142 -54
rect 154 -58 158 -54
rect 212 -68 216 -64
rect 220 -68 224 -64
rect 252 -68 256 -64
rect 260 -68 264 -64
rect 268 -68 272 -64
rect 276 -68 280 -64
rect 51 -72 55 -68
rect 62 -72 66 -68
rect 72 -72 76 -68
rect -13 -208 -9 -204
rect -3 -208 1 -204
rect 7 -208 11 -204
rect 58 -225 62 -221
rect 69 -225 73 -221
rect 79 -225 83 -221
rect 90 -225 94 -221
rect 132 -242 136 -238
rect 142 -242 146 -238
rect 154 -242 158 -238
rect 166 -242 170 -238
rect 176 -242 180 -238
rect 240 -259 244 -255
rect 250 -259 254 -255
rect 262 -259 266 -255
rect 274 -259 278 -255
rect 286 -259 290 -255
rect 296 -259 300 -255
rect 150 -328 154 -324
rect 158 -328 162 -324
rect 190 -328 194 -324
rect 198 -328 202 -324
rect 206 -328 210 -324
rect 214 -328 218 -324
rect -13 -391 -9 -387
rect -5 -391 -1 -387
rect 27 -391 31 -387
rect 35 -391 39 -387
rect 43 -391 47 -387
rect 51 -391 55 -387
rect 66 -408 70 -404
rect 76 -408 80 -404
rect 86 -408 90 -404
rect 101 -408 105 -404
rect 111 -408 115 -404
rect 121 -408 125 -404
rect 169 -423 173 -419
rect 177 -423 181 -419
rect 209 -423 213 -419
rect 217 -423 221 -419
rect 225 -423 229 -419
rect 233 -423 237 -419
rect 15 -461 19 -457
rect 25 -461 29 -457
rect -13 -478 -9 -474
rect -3 -478 1 -474
rect 7 -478 11 -474
rect 75 -572 79 -568
rect 85 -572 89 -568
rect 97 -572 101 -568
rect 107 -572 111 -568
rect 129 -572 133 -568
rect 139 -572 143 -568
rect 151 -572 155 -568
rect 161 -572 165 -568
rect -13 -580 -9 -576
rect -5 -580 -1 -576
rect 27 -580 31 -576
rect 35 -580 39 -576
rect 43 -580 47 -576
rect 15 -650 19 -646
rect 25 -650 29 -646
rect 151 -650 155 -646
rect 159 -650 163 -646
rect 191 -650 195 -646
rect 199 -650 203 -646
rect 207 -650 211 -646
rect 215 -650 219 -646
rect 75 -659 79 -655
rect 85 -659 89 -655
rect 95 -659 99 -655
rect -13 -667 -9 -663
rect -3 -667 1 -663
rect 7 -667 11 -663
rect 81 -789 85 -785
rect 91 -789 95 -785
rect 103 -789 107 -785
rect 115 -789 119 -785
rect 125 -789 129 -785
rect -13 -816 -9 -812
rect -5 -816 -1 -812
rect 27 -816 31 -812
rect 35 -816 39 -812
rect 43 -816 47 -812
rect 51 -816 55 -812
rect 221 -816 225 -812
rect 229 -816 233 -812
rect 261 -816 265 -812
rect 269 -816 273 -812
rect 277 -816 281 -812
rect 285 -816 289 -812
rect 151 -853 155 -849
rect 161 -853 165 -849
rect 173 -853 177 -849
rect 185 -853 189 -849
rect 195 -853 199 -849
rect 15 -886 19 -882
rect 25 -886 29 -882
rect 87 -893 91 -889
rect 98 -893 102 -889
rect 108 -893 112 -889
rect 119 -893 123 -889
rect -13 -903 -9 -899
rect -3 -903 1 -899
rect 7 -903 11 -899
rect 87 -980 91 -976
rect 97 -980 101 -976
rect 107 -980 111 -976
rect 75 -1126 79 -1122
rect 85 -1126 89 -1122
rect 97 -1126 101 -1122
rect 109 -1126 113 -1122
rect 121 -1126 125 -1122
rect 131 -1126 135 -1122
rect -13 -1197 -9 -1193
rect -5 -1197 -1 -1193
rect 27 -1197 31 -1193
rect 35 -1197 39 -1193
rect 43 -1197 47 -1193
rect 51 -1197 55 -1193
rect 83 -1249 87 -1245
rect 93 -1249 97 -1245
rect 105 -1249 109 -1245
rect 117 -1249 121 -1245
rect 127 -1249 131 -1245
rect 15 -1267 19 -1263
rect 25 -1267 29 -1263
rect 154 -1266 158 -1262
rect 164 -1266 168 -1262
rect 176 -1266 180 -1262
rect 188 -1266 192 -1262
rect 200 -1266 204 -1262
rect 210 -1266 214 -1262
rect -13 -1284 -9 -1280
rect -3 -1284 1 -1280
rect 7 -1284 11 -1280
rect 93 -1355 97 -1351
rect 104 -1355 108 -1351
rect 114 -1355 118 -1351
rect 125 -1355 129 -1351
rect 103 -1443 107 -1439
rect 113 -1443 117 -1439
rect 123 -1443 127 -1439
<< nsubstratencontact >>
rect 53 16 57 20
rect 65 16 69 20
rect 76 16 80 20
rect 87 16 91 20
rect 101 16 105 20
rect 112 16 116 20
rect 122 16 126 20
rect 136 16 140 20
rect 152 16 156 20
rect 164 16 168 20
rect -20 7 -16 11
rect -12 7 -8 11
rect 252 -8 256 -4
rect 268 -8 272 -4
rect -13 -131 -9 -127
rect -3 -131 1 -127
rect 7 -131 11 -127
rect 58 -131 62 -127
rect 69 -131 73 -127
rect 80 -131 84 -127
rect 90 -131 94 -127
rect 132 -131 136 -127
rect 143 -131 147 -127
rect 154 -131 158 -127
rect 165 -131 169 -127
rect 176 -131 180 -127
rect 240 -131 244 -127
rect 251 -131 255 -127
rect 262 -131 266 -127
rect 273 -131 277 -127
rect 286 -131 290 -127
rect 296 -131 300 -127
rect 27 -331 31 -327
rect 43 -331 47 -327
rect 66 -331 70 -327
rect 76 -331 80 -327
rect 86 -331 90 -327
rect 101 -331 105 -327
rect 111 -331 115 -327
rect 121 -331 125 -327
rect -13 -401 -9 -397
rect -3 -401 1 -397
rect 7 -401 11 -397
rect 15 -401 19 -397
rect 25 -401 29 -397
rect 190 -388 194 -384
rect 206 -388 210 -384
rect 75 -478 79 -474
rect 86 -478 90 -474
rect 97 -478 101 -474
rect 107 -478 111 -474
rect 129 -478 133 -474
rect 140 -478 144 -474
rect 151 -478 155 -474
rect 161 -478 165 -474
rect 209 -483 213 -479
rect 225 -483 229 -479
rect 27 -520 31 -516
rect 43 -520 47 -516
rect 75 -582 79 -578
rect 85 -582 89 -578
rect 95 -582 99 -578
rect -13 -590 -9 -586
rect -3 -590 1 -586
rect 7 -590 11 -586
rect 15 -590 19 -586
rect 23 -590 27 -586
rect 81 -678 85 -674
rect 92 -678 96 -674
rect 103 -678 107 -674
rect 114 -678 118 -674
rect 125 -678 129 -674
rect 191 -710 195 -706
rect 207 -710 211 -706
rect 27 -756 31 -752
rect 43 -756 47 -752
rect 151 -742 155 -738
rect 162 -742 166 -738
rect 173 -742 177 -738
rect 184 -742 188 -738
rect 195 -742 199 -738
rect 87 -799 91 -795
rect 98 -799 102 -795
rect 109 -799 113 -795
rect 119 -799 123 -795
rect 261 -756 265 -752
rect 277 -756 281 -752
rect -13 -826 -9 -822
rect -3 -826 1 -822
rect 7 -826 11 -822
rect 15 -826 19 -822
rect 25 -826 29 -822
rect 87 -903 91 -899
rect 97 -903 101 -899
rect 107 -903 111 -899
rect 75 -998 79 -994
rect 86 -998 90 -994
rect 97 -998 101 -994
rect 108 -998 112 -994
rect 121 -998 125 -994
rect 131 -998 135 -994
rect 27 -1137 31 -1133
rect 43 -1137 47 -1133
rect 83 -1138 87 -1134
rect 94 -1138 98 -1134
rect 105 -1138 109 -1134
rect 116 -1138 120 -1134
rect 127 -1138 131 -1134
rect 154 -1138 158 -1134
rect 165 -1138 169 -1134
rect 176 -1138 180 -1134
rect 187 -1138 191 -1134
rect 200 -1138 204 -1134
rect 210 -1138 214 -1134
rect -13 -1207 -9 -1203
rect -3 -1207 1 -1203
rect 7 -1207 11 -1203
rect 15 -1207 19 -1203
rect 25 -1207 29 -1203
rect 93 -1261 97 -1257
rect 104 -1261 108 -1257
rect 115 -1261 119 -1257
rect 125 -1261 129 -1257
rect 103 -1366 107 -1362
rect 113 -1366 117 -1362
rect 123 -1366 127 -1362
<< polysilicon >>
rect 60 10 62 13
rect 72 10 74 13
rect 96 10 98 13
rect 131 10 133 13
rect 159 10 161 13
rect 217 11 219 14
rect 233 11 235 14
rect -15 1 -13 4
rect -15 -35 -13 -19
rect 96 -30 98 -10
rect 108 -30 110 -23
rect 131 -30 133 -10
rect 143 -30 145 -23
rect 159 -26 161 -10
rect -15 -48 -13 -45
rect 60 -54 62 -30
rect 72 -44 74 -30
rect 257 -14 259 -11
rect 273 -14 275 -11
rect 159 -39 161 -36
rect 217 -50 219 -29
rect 233 -40 235 -29
rect 257 -50 259 -34
rect 273 -50 275 -34
rect 96 -53 98 -50
rect 108 -53 110 -50
rect 131 -53 133 -50
rect 143 -53 145 -50
rect 217 -63 219 -60
rect 257 -63 259 -60
rect 273 -63 275 -60
rect 60 -67 62 -64
rect -8 -137 -6 -134
rect 4 -137 6 -134
rect 63 -137 65 -134
rect 75 -137 77 -134
rect 87 -137 89 -134
rect 137 -137 139 -134
rect 149 -137 151 -134
rect 161 -137 163 -134
rect 173 -137 175 -134
rect 245 -137 247 -134
rect 257 -137 259 -134
rect 269 -137 271 -134
rect 281 -137 283 -134
rect 293 -137 295 -134
rect -8 -180 -6 -157
rect 4 -180 6 -157
rect 63 -187 65 -157
rect 75 -187 77 -157
rect 87 -187 89 -157
rect -8 -203 -6 -200
rect 4 -203 6 -200
rect 137 -194 139 -157
rect 149 -194 151 -157
rect 161 -194 163 -157
rect 173 -194 175 -157
rect 63 -220 65 -217
rect 75 -220 77 -217
rect 87 -220 89 -217
rect 245 -201 247 -157
rect 257 -201 259 -157
rect 269 -201 271 -157
rect 281 -201 283 -157
rect 293 -201 295 -157
rect 137 -237 139 -234
rect 149 -237 151 -234
rect 161 -237 163 -234
rect 173 -237 175 -234
rect 245 -254 247 -251
rect 257 -254 259 -251
rect 269 -254 271 -251
rect 281 -254 283 -251
rect 293 -254 295 -251
rect -8 -312 -6 -309
rect 8 -312 10 -309
rect 155 -332 157 -329
rect 195 -332 197 -329
rect 211 -332 213 -329
rect 32 -337 34 -334
rect 48 -337 50 -334
rect 71 -337 73 -334
rect 83 -337 85 -334
rect 106 -337 108 -334
rect 118 -337 120 -334
rect -8 -373 -6 -352
rect 8 -363 10 -352
rect 32 -373 34 -357
rect 48 -373 50 -357
rect 71 -380 73 -357
rect 83 -380 85 -357
rect 106 -380 108 -357
rect 118 -380 120 -357
rect 155 -363 157 -342
rect 171 -363 173 -352
rect 195 -358 197 -342
rect 211 -358 213 -342
rect -8 -386 -6 -383
rect 32 -386 34 -383
rect 48 -386 50 -383
rect 71 -403 73 -400
rect 83 -403 85 -400
rect 106 -403 108 -400
rect 118 -403 120 -400
rect 195 -381 197 -378
rect 211 -381 213 -378
rect -8 -407 -6 -404
rect 4 -407 6 -404
rect 20 -407 22 -404
rect 155 -406 157 -403
rect 171 -406 173 -403
rect 174 -427 176 -424
rect 214 -427 216 -424
rect 230 -427 232 -424
rect -8 -450 -6 -427
rect 4 -450 6 -427
rect 20 -443 22 -427
rect 20 -456 22 -453
rect 174 -458 176 -437
rect 190 -458 192 -447
rect 214 -453 216 -437
rect 230 -453 232 -437
rect -8 -473 -6 -470
rect 4 -473 6 -470
rect 80 -484 82 -481
rect 92 -484 94 -481
rect 104 -484 106 -481
rect 134 -484 136 -481
rect 146 -484 148 -481
rect 158 -484 160 -481
rect -8 -501 -6 -498
rect 8 -501 10 -498
rect 214 -476 216 -473
rect 230 -476 232 -473
rect 174 -501 176 -498
rect 190 -501 192 -498
rect 32 -526 34 -523
rect 48 -526 50 -523
rect -8 -562 -6 -541
rect 8 -552 10 -541
rect 80 -534 82 -504
rect 92 -534 94 -504
rect 104 -534 106 -504
rect 134 -534 136 -504
rect 146 -534 148 -504
rect 158 -534 160 -504
rect 32 -562 34 -546
rect 48 -562 50 -546
rect 80 -567 82 -564
rect 92 -567 94 -564
rect 104 -567 106 -564
rect 134 -567 136 -564
rect 146 -567 148 -564
rect 158 -567 160 -564
rect -8 -575 -6 -572
rect 32 -575 34 -572
rect 48 -575 50 -572
rect 80 -588 82 -585
rect 92 -588 94 -585
rect -8 -596 -6 -593
rect 4 -596 6 -593
rect 20 -596 22 -593
rect -8 -639 -6 -616
rect 4 -639 6 -616
rect 20 -632 22 -616
rect 80 -631 82 -608
rect 92 -631 94 -608
rect 20 -645 22 -642
rect 80 -654 82 -651
rect 92 -654 94 -651
rect 156 -654 158 -651
rect 196 -654 198 -651
rect 212 -654 214 -651
rect -8 -662 -6 -659
rect 4 -662 6 -659
rect 86 -684 88 -681
rect 98 -684 100 -681
rect 110 -684 112 -681
rect 122 -684 124 -681
rect 156 -685 158 -664
rect 172 -685 174 -674
rect 196 -680 198 -664
rect 212 -680 214 -664
rect -8 -737 -6 -734
rect 8 -737 10 -734
rect 86 -741 88 -704
rect 98 -741 100 -704
rect 110 -741 112 -704
rect 122 -741 124 -704
rect 196 -703 198 -700
rect 212 -703 214 -700
rect 156 -728 158 -725
rect 172 -728 174 -725
rect 226 -737 228 -734
rect 242 -737 244 -734
rect 32 -762 34 -759
rect 48 -762 50 -759
rect -8 -798 -6 -777
rect 8 -788 10 -777
rect 156 -748 158 -745
rect 168 -748 170 -745
rect 180 -748 182 -745
rect 192 -748 194 -745
rect 32 -798 34 -782
rect 48 -798 50 -782
rect 86 -784 88 -781
rect 98 -784 100 -781
rect 110 -784 112 -781
rect 122 -784 124 -781
rect 92 -805 94 -802
rect 104 -805 106 -802
rect 116 -805 118 -802
rect 156 -805 158 -768
rect 168 -805 170 -768
rect 180 -805 182 -768
rect 192 -805 194 -768
rect 266 -762 268 -759
rect 282 -762 284 -759
rect 226 -798 228 -777
rect 242 -788 244 -777
rect 266 -798 268 -782
rect 282 -798 284 -782
rect -8 -811 -6 -808
rect 32 -811 34 -808
rect 48 -811 50 -808
rect -8 -832 -6 -829
rect 4 -832 6 -829
rect 20 -832 22 -829
rect -8 -875 -6 -852
rect 4 -875 6 -852
rect 20 -868 22 -852
rect 92 -855 94 -825
rect 104 -855 106 -825
rect 116 -855 118 -825
rect 226 -811 228 -808
rect 266 -811 268 -808
rect 282 -811 284 -808
rect 156 -848 158 -845
rect 168 -848 170 -845
rect 180 -848 182 -845
rect 192 -848 194 -845
rect 20 -881 22 -878
rect 92 -888 94 -885
rect 104 -888 106 -885
rect 116 -888 118 -885
rect -8 -898 -6 -895
rect 4 -898 6 -895
rect 92 -909 94 -906
rect 104 -909 106 -906
rect 92 -952 94 -929
rect 104 -952 106 -929
rect 92 -975 94 -972
rect 104 -975 106 -972
rect 80 -1004 82 -1001
rect 92 -1004 94 -1001
rect 104 -1004 106 -1001
rect 116 -1004 118 -1001
rect 128 -1004 130 -1001
rect 80 -1068 82 -1024
rect 92 -1068 94 -1024
rect 104 -1068 106 -1024
rect 116 -1068 118 -1024
rect 128 -1068 130 -1024
rect -8 -1118 -6 -1115
rect 8 -1118 10 -1115
rect 80 -1121 82 -1118
rect 92 -1121 94 -1118
rect 104 -1121 106 -1118
rect 116 -1121 118 -1118
rect 128 -1121 130 -1118
rect 32 -1143 34 -1140
rect 48 -1143 50 -1140
rect -8 -1179 -6 -1158
rect 8 -1169 10 -1158
rect 88 -1144 90 -1141
rect 100 -1144 102 -1141
rect 112 -1144 114 -1141
rect 124 -1144 126 -1141
rect 159 -1144 161 -1141
rect 171 -1144 173 -1141
rect 183 -1144 185 -1141
rect 195 -1144 197 -1141
rect 207 -1144 209 -1141
rect 32 -1179 34 -1163
rect 48 -1179 50 -1163
rect -8 -1192 -6 -1189
rect 32 -1192 34 -1189
rect 48 -1192 50 -1189
rect 88 -1201 90 -1164
rect 100 -1201 102 -1164
rect 112 -1201 114 -1164
rect 124 -1201 126 -1164
rect -8 -1213 -6 -1210
rect 4 -1213 6 -1210
rect 20 -1213 22 -1210
rect -8 -1256 -6 -1233
rect 4 -1256 6 -1233
rect 20 -1249 22 -1233
rect 159 -1208 161 -1164
rect 171 -1208 173 -1164
rect 183 -1208 185 -1164
rect 195 -1208 197 -1164
rect 207 -1208 209 -1164
rect 88 -1244 90 -1241
rect 100 -1244 102 -1241
rect 112 -1244 114 -1241
rect 124 -1244 126 -1241
rect 20 -1262 22 -1259
rect 159 -1261 161 -1258
rect 171 -1261 173 -1258
rect 183 -1261 185 -1258
rect 195 -1261 197 -1258
rect 207 -1261 209 -1258
rect 98 -1267 100 -1264
rect 110 -1267 112 -1264
rect 122 -1267 124 -1264
rect -8 -1279 -6 -1276
rect 4 -1279 6 -1276
rect 98 -1317 100 -1287
rect 110 -1317 112 -1287
rect 122 -1317 124 -1287
rect 98 -1350 100 -1347
rect 110 -1350 112 -1347
rect 122 -1350 124 -1347
rect 108 -1372 110 -1369
rect 120 -1372 122 -1369
rect 108 -1415 110 -1392
rect 120 -1415 122 -1392
rect 108 -1438 110 -1435
rect 120 -1438 122 -1435
<< polycontact >>
rect -19 -32 -15 -28
rect 92 -20 96 -16
rect 127 -21 131 -17
rect 104 -27 108 -23
rect 155 -23 159 -19
rect 139 -27 143 -23
rect 56 -51 60 -47
rect 68 -42 72 -38
rect 213 -47 217 -43
rect 229 -40 233 -36
rect 253 -47 257 -43
rect 269 -47 273 -43
rect -12 -170 -8 -166
rect 0 -177 4 -173
rect 59 -170 63 -166
rect 71 -177 75 -173
rect 83 -184 87 -180
rect 133 -170 137 -166
rect 145 -177 149 -173
rect 157 -184 161 -180
rect 169 -191 173 -187
rect 241 -170 245 -166
rect 253 -177 257 -173
rect 265 -184 269 -180
rect 277 -191 281 -187
rect 289 -198 293 -194
rect -12 -370 -8 -366
rect 4 -363 8 -359
rect 151 -349 155 -345
rect 28 -370 32 -366
rect 44 -370 48 -366
rect 67 -370 71 -366
rect 79 -377 83 -373
rect 102 -370 106 -366
rect 114 -377 118 -373
rect 191 -349 195 -345
rect 167 -356 171 -352
rect 207 -349 211 -345
rect -12 -440 -8 -436
rect 0 -447 4 -443
rect 16 -440 20 -436
rect 170 -444 174 -440
rect 210 -444 214 -440
rect 186 -451 190 -447
rect 226 -444 230 -440
rect 76 -517 80 -513
rect -12 -559 -8 -555
rect 4 -552 8 -548
rect 88 -524 92 -520
rect 100 -531 104 -527
rect 130 -517 134 -513
rect 142 -524 146 -520
rect 154 -531 158 -527
rect 28 -559 32 -555
rect 44 -559 48 -555
rect -12 -629 -8 -625
rect 0 -636 4 -632
rect 16 -629 20 -625
rect 76 -621 80 -617
rect 88 -628 92 -624
rect 152 -671 156 -667
rect 192 -671 196 -667
rect 168 -678 172 -674
rect 208 -671 212 -667
rect 82 -717 86 -713
rect 94 -724 98 -720
rect 106 -731 110 -727
rect 118 -738 122 -734
rect -12 -795 -8 -791
rect 4 -788 8 -784
rect 152 -781 156 -777
rect 28 -795 32 -791
rect 44 -795 48 -791
rect 164 -788 168 -784
rect 176 -795 180 -791
rect 188 -802 192 -798
rect 222 -795 226 -791
rect 238 -788 242 -784
rect 262 -795 266 -791
rect 278 -795 282 -791
rect 88 -838 92 -834
rect -12 -865 -8 -861
rect 0 -872 4 -868
rect 16 -865 20 -861
rect 100 -845 104 -841
rect 112 -852 116 -848
rect 88 -942 92 -938
rect 100 -949 104 -945
rect 76 -1037 80 -1033
rect 88 -1044 92 -1040
rect 100 -1051 104 -1047
rect 112 -1058 116 -1054
rect 124 -1065 128 -1061
rect -12 -1176 -8 -1172
rect 4 -1169 8 -1165
rect 28 -1176 32 -1172
rect 44 -1176 48 -1172
rect 84 -1177 88 -1173
rect 96 -1184 100 -1180
rect 108 -1191 112 -1187
rect 120 -1198 124 -1194
rect 155 -1177 159 -1173
rect -12 -1246 -8 -1242
rect 0 -1253 4 -1249
rect 16 -1246 20 -1242
rect 167 -1184 171 -1180
rect 179 -1191 183 -1187
rect 191 -1198 195 -1194
rect 203 -1205 207 -1201
rect 94 -1300 98 -1296
rect 106 -1307 110 -1303
rect 118 -1314 122 -1310
rect 104 -1405 108 -1401
rect 116 -1412 120 -1408
<< metal1 >>
rect 49 16 53 20
rect 57 16 65 20
rect 69 16 76 20
rect 80 16 87 20
rect 91 16 101 20
rect 105 16 112 20
rect 116 16 122 20
rect 126 16 136 20
rect 140 16 152 20
rect 156 16 164 20
rect 168 16 172 20
rect 212 17 246 21
rect -16 7 -12 11
rect 55 10 59 16
rect 91 10 95 16
rect 126 10 130 16
rect 154 10 158 16
rect 212 11 216 17
rect 228 11 232 17
rect -20 1 -16 7
rect -12 -28 -8 -19
rect -26 -32 -19 -28
rect -12 -32 -2 -28
rect 90 -20 92 -16
rect 99 -17 103 -10
rect 134 -17 138 -10
rect 99 -20 127 -17
rect 111 -21 127 -20
rect 134 -19 150 -17
rect 162 -19 166 -10
rect 134 -20 155 -19
rect 79 -27 104 -24
rect 111 -30 115 -21
rect 146 -23 155 -20
rect 162 -23 172 -19
rect 123 -27 139 -24
rect 146 -30 150 -23
rect 162 -26 166 -23
rect -12 -35 -8 -32
rect 49 -42 53 -38
rect 58 -42 68 -38
rect -20 -49 -16 -45
rect 75 -47 79 -30
rect -16 -53 -12 -49
rect 49 -51 56 -47
rect 63 -51 79 -47
rect 221 -36 224 -29
rect 154 -40 158 -36
rect 206 -40 229 -36
rect 158 -44 164 -40
rect 168 -44 172 -40
rect 237 -43 240 -29
rect 63 -54 67 -51
rect 91 -54 95 -50
rect 126 -54 130 -50
rect 154 -54 158 -44
rect 206 -47 213 -43
rect 217 -47 240 -43
rect 243 -43 246 17
rect 256 -8 268 -4
rect 252 -14 256 -8
rect 268 -14 272 -8
rect 260 -43 264 -34
rect 276 -43 280 -34
rect 243 -47 253 -43
rect 260 -47 269 -43
rect 276 -47 286 -43
rect 243 -50 246 -47
rect 260 -50 264 -47
rect 276 -50 280 -47
rect 76 -58 87 -54
rect 91 -58 103 -54
rect 107 -58 122 -54
rect 126 -58 138 -54
rect 142 -58 154 -54
rect 55 -68 59 -64
rect 72 -68 76 -58
rect 224 -53 246 -50
rect 212 -64 216 -60
rect 252 -64 256 -60
rect 268 -64 272 -60
rect 216 -68 220 -64
rect 224 -68 252 -64
rect 256 -68 260 -64
rect 264 -68 268 -64
rect 272 -68 276 -64
rect 49 -72 51 -68
rect 55 -72 62 -68
rect 66 -72 72 -68
rect -9 -131 -3 -127
rect 1 -131 7 -127
rect -13 -137 -9 -131
rect 7 -137 11 -131
rect 62 -131 69 -127
rect 73 -131 80 -127
rect 84 -131 90 -127
rect 136 -131 143 -127
rect 147 -131 154 -127
rect 158 -131 165 -127
rect 169 -131 176 -127
rect 58 -137 62 -131
rect 80 -137 84 -131
rect 132 -137 136 -131
rect 154 -137 158 -131
rect 176 -137 180 -131
rect 244 -131 251 -127
rect 255 -131 262 -127
rect 266 -131 273 -127
rect 277 -131 286 -127
rect 290 -131 296 -127
rect 240 -137 244 -131
rect 262 -137 266 -131
rect 286 -137 290 -131
rect -3 -166 1 -157
rect 68 -166 72 -157
rect 90 -166 94 -157
rect 142 -160 146 -157
rect 166 -160 170 -157
rect 142 -163 170 -160
rect 250 -160 254 -157
rect 274 -160 278 -157
rect 296 -160 300 -157
rect 250 -163 300 -160
rect -19 -170 -12 -166
rect -3 -170 17 -166
rect 52 -170 59 -166
rect 68 -170 94 -166
rect 126 -170 133 -166
rect -19 -177 0 -173
rect 7 -180 11 -170
rect 90 -173 94 -170
rect 166 -173 170 -163
rect 234 -170 241 -166
rect 52 -177 71 -173
rect 90 -177 100 -173
rect 126 -177 145 -173
rect 166 -177 186 -173
rect 234 -177 253 -173
rect 52 -184 83 -180
rect 90 -187 94 -177
rect 126 -184 157 -180
rect -13 -204 -9 -200
rect -9 -208 -3 -204
rect 1 -208 7 -204
rect 126 -191 169 -187
rect 176 -194 180 -177
rect 296 -180 300 -163
rect 234 -184 265 -180
rect 296 -184 306 -180
rect 234 -191 277 -187
rect 58 -221 62 -217
rect 62 -225 69 -221
rect 73 -225 79 -221
rect 83 -225 90 -221
rect 234 -198 289 -194
rect 296 -201 300 -184
rect 132 -238 136 -234
rect 136 -242 142 -238
rect 146 -242 154 -238
rect 158 -242 166 -238
rect 170 -242 176 -238
rect 240 -255 244 -251
rect 244 -259 250 -255
rect 254 -259 262 -255
rect 266 -259 274 -255
rect 278 -259 286 -255
rect 290 -259 296 -255
rect -13 -306 21 -302
rect -13 -312 -9 -306
rect 3 -312 7 -306
rect -4 -359 -1 -352
rect -27 -362 4 -359
rect -27 -436 -24 -362
rect 12 -366 15 -352
rect -16 -370 -12 -366
rect -8 -370 15 -366
rect 18 -366 21 -306
rect 31 -331 43 -327
rect 27 -337 31 -331
rect 43 -337 47 -331
rect 70 -331 76 -327
rect 80 -331 86 -327
rect 90 -330 101 -327
rect 66 -337 70 -331
rect 86 -337 90 -331
rect 105 -331 111 -327
rect 115 -331 121 -327
rect 101 -337 105 -331
rect 121 -337 125 -331
rect 154 -328 158 -324
rect 162 -328 190 -324
rect 194 -328 198 -324
rect 202 -328 206 -324
rect 210 -328 214 -324
rect 150 -332 154 -328
rect 190 -332 194 -328
rect 206 -332 210 -328
rect 162 -342 184 -339
rect 181 -345 184 -342
rect 198 -345 202 -342
rect 214 -345 218 -342
rect 137 -349 151 -345
rect 155 -349 178 -345
rect 144 -356 167 -352
rect 35 -366 39 -357
rect 51 -366 55 -357
rect 18 -370 28 -366
rect 35 -370 44 -366
rect 51 -370 58 -366
rect 76 -366 80 -357
rect 111 -366 115 -357
rect 63 -370 67 -366
rect 76 -370 102 -366
rect 111 -370 125 -366
rect 18 -373 21 -370
rect 35 -373 39 -370
rect 51 -373 55 -370
rect -1 -376 21 -373
rect 60 -377 79 -373
rect -13 -387 -9 -383
rect 27 -387 31 -383
rect 43 -387 47 -383
rect -9 -391 -5 -387
rect -1 -391 27 -387
rect 31 -391 35 -387
rect 39 -391 43 -387
rect 47 -391 51 -387
rect -9 -401 -3 -397
rect 1 -401 7 -397
rect 11 -401 15 -397
rect 19 -401 25 -397
rect 29 -401 33 -397
rect -13 -407 -9 -401
rect 7 -407 11 -401
rect 15 -407 19 -401
rect -3 -436 1 -427
rect 23 -436 27 -427
rect 60 -411 63 -377
rect 86 -380 90 -370
rect 98 -377 114 -373
rect 121 -380 125 -370
rect 125 -400 128 -397
rect 66 -404 70 -400
rect 101 -404 105 -400
rect 70 -408 76 -404
rect 80 -408 86 -404
rect 90 -408 101 -404
rect 105 -408 111 -404
rect 115 -408 121 -404
rect 144 -411 147 -356
rect 159 -363 162 -356
rect 175 -363 178 -349
rect 60 -414 147 -411
rect 181 -349 191 -345
rect 198 -349 207 -345
rect 214 -349 224 -345
rect 150 -409 154 -403
rect 166 -409 170 -403
rect 181 -409 184 -349
rect 198 -358 202 -349
rect 214 -358 218 -349
rect 190 -384 194 -378
rect 206 -384 210 -378
rect 194 -388 206 -384
rect 150 -413 184 -409
rect -27 -439 -12 -436
rect -3 -440 16 -436
rect 23 -439 41 -436
rect -16 -447 0 -444
rect 7 -450 11 -440
rect 23 -443 27 -439
rect 15 -457 19 -453
rect 19 -461 25 -457
rect 11 -470 30 -466
rect -13 -474 -9 -470
rect -9 -478 -3 -474
rect 1 -478 7 -474
rect -13 -495 21 -491
rect 38 -494 41 -439
rect -13 -501 -9 -495
rect 3 -501 7 -495
rect -4 -548 -1 -541
rect -27 -551 4 -548
rect -27 -625 -24 -551
rect 12 -555 15 -541
rect -16 -559 -12 -555
rect -8 -559 15 -555
rect 18 -555 21 -495
rect 31 -520 43 -516
rect 27 -526 31 -520
rect 43 -526 47 -520
rect 51 -526 54 -452
rect 60 -512 63 -414
rect 173 -423 177 -419
rect 181 -423 209 -419
rect 213 -423 217 -419
rect 221 -423 225 -419
rect 229 -423 233 -419
rect 169 -427 173 -423
rect 209 -427 213 -423
rect 225 -427 229 -423
rect 181 -437 203 -434
rect 200 -440 203 -437
rect 217 -440 221 -437
rect 233 -440 237 -437
rect 134 -444 170 -441
rect 174 -444 197 -440
rect 163 -448 186 -447
rect 155 -451 186 -448
rect 178 -458 181 -451
rect 194 -458 197 -444
rect 79 -478 86 -474
rect 90 -478 97 -474
rect 101 -478 107 -474
rect 111 -478 129 -474
rect 133 -478 140 -474
rect 144 -478 151 -474
rect 155 -478 161 -474
rect 75 -484 79 -478
rect 97 -484 101 -478
rect 129 -484 133 -478
rect 151 -484 155 -478
rect 85 -513 89 -504
rect 107 -513 111 -504
rect 139 -513 143 -504
rect 161 -513 165 -504
rect 200 -444 210 -440
rect 217 -444 226 -440
rect 233 -444 243 -440
rect 169 -504 173 -498
rect 185 -504 189 -498
rect 200 -504 203 -444
rect 217 -453 221 -444
rect 233 -453 237 -444
rect 209 -479 213 -473
rect 225 -479 229 -473
rect 213 -483 225 -479
rect 169 -508 203 -504
rect 65 -517 76 -513
rect 85 -517 130 -513
rect 139 -517 165 -513
rect 87 -524 88 -520
rect 35 -555 39 -546
rect 51 -555 55 -546
rect 63 -531 100 -528
rect 63 -555 66 -531
rect 107 -534 111 -517
rect 18 -559 28 -555
rect 35 -559 44 -555
rect 51 -558 66 -555
rect 18 -562 21 -559
rect 35 -562 39 -559
rect 51 -562 55 -558
rect -1 -565 21 -562
rect -13 -576 -9 -572
rect 27 -576 31 -572
rect 43 -576 47 -572
rect 61 -559 66 -558
rect 51 -576 54 -572
rect -9 -580 -5 -576
rect -1 -580 27 -576
rect 31 -580 35 -576
rect 39 -580 43 -576
rect -9 -590 -3 -586
rect 1 -590 7 -586
rect 11 -590 15 -586
rect 19 -590 23 -586
rect -13 -596 -9 -590
rect 7 -596 11 -590
rect 15 -596 19 -590
rect -3 -625 1 -616
rect 23 -625 27 -616
rect 61 -624 64 -559
rect 115 -524 142 -520
rect 75 -568 79 -564
rect 79 -572 85 -568
rect 89 -572 97 -568
rect 101 -572 107 -568
rect 79 -582 85 -578
rect 89 -582 95 -578
rect 75 -588 79 -582
rect 95 -588 99 -582
rect 72 -617 75 -611
rect 85 -617 89 -608
rect 115 -617 118 -524
rect 72 -621 76 -617
rect 85 -621 118 -617
rect 122 -531 154 -527
rect -27 -628 -12 -625
rect -3 -629 16 -625
rect -16 -636 0 -633
rect 7 -639 11 -629
rect 61 -628 88 -624
rect 23 -632 27 -630
rect 95 -631 99 -621
rect 15 -646 19 -642
rect 19 -650 25 -646
rect 75 -655 79 -651
rect 11 -659 34 -656
rect 79 -659 85 -655
rect 89 -659 95 -655
rect -13 -663 -9 -659
rect 31 -662 34 -659
rect 122 -662 125 -531
rect 161 -534 165 -517
rect 165 -564 171 -561
rect 129 -568 133 -564
rect 133 -572 139 -568
rect 143 -572 151 -568
rect 155 -572 161 -568
rect 168 -575 171 -564
rect -9 -667 -3 -663
rect 1 -667 7 -663
rect 31 -665 125 -662
rect 145 -578 171 -575
rect 145 -667 148 -578
rect 155 -650 159 -646
rect 163 -650 191 -646
rect 195 -650 199 -646
rect 203 -650 207 -646
rect 211 -650 215 -646
rect 151 -654 155 -650
rect 191 -654 195 -650
rect 207 -654 211 -650
rect 163 -664 185 -661
rect 182 -667 185 -664
rect 199 -667 203 -664
rect 215 -667 219 -664
rect 74 -671 138 -668
rect 145 -671 152 -667
rect 156 -671 179 -667
rect 74 -713 77 -671
rect 135 -674 138 -671
rect 85 -678 92 -674
rect 96 -678 103 -674
rect 107 -678 114 -674
rect 118 -678 125 -674
rect 135 -678 168 -674
rect 81 -684 85 -678
rect 103 -684 107 -678
rect 125 -684 129 -678
rect 160 -685 163 -678
rect 176 -685 179 -671
rect 91 -707 95 -704
rect 115 -707 119 -704
rect 91 -710 119 -707
rect 52 -716 82 -713
rect -13 -731 21 -727
rect -13 -737 -9 -731
rect 3 -737 7 -731
rect -4 -784 -1 -777
rect -27 -787 4 -784
rect -27 -861 -24 -787
rect 12 -791 15 -777
rect -16 -795 -12 -791
rect -8 -795 15 -791
rect 18 -791 21 -731
rect 31 -756 43 -752
rect 27 -762 31 -756
rect 43 -762 47 -756
rect 52 -762 55 -716
rect 115 -720 119 -710
rect 79 -724 94 -720
rect 115 -724 129 -720
rect 63 -731 106 -728
rect 72 -738 118 -735
rect 35 -791 39 -782
rect 51 -791 55 -782
rect 18 -795 28 -791
rect 35 -795 44 -791
rect 51 -795 61 -791
rect 18 -798 21 -795
rect 35 -798 39 -795
rect 51 -798 55 -795
rect -1 -801 21 -798
rect -13 -812 -9 -808
rect 27 -812 31 -808
rect 43 -812 47 -808
rect -9 -816 -5 -812
rect -1 -816 27 -812
rect 31 -816 35 -812
rect 39 -816 43 -812
rect 47 -816 51 -812
rect -9 -826 -3 -822
rect 1 -826 7 -822
rect 11 -826 15 -822
rect 19 -826 25 -822
rect 29 -826 33 -822
rect -13 -832 -9 -826
rect 7 -832 11 -826
rect 15 -832 19 -826
rect 58 -848 61 -795
rect 75 -833 78 -738
rect 125 -741 129 -724
rect 182 -671 192 -667
rect 199 -671 208 -667
rect 215 -671 225 -667
rect 151 -731 155 -725
rect 167 -731 171 -725
rect 182 -731 185 -671
rect 199 -680 203 -671
rect 215 -680 219 -671
rect 191 -706 195 -700
rect 207 -706 211 -700
rect 195 -710 207 -706
rect 151 -735 185 -731
rect 221 -731 255 -727
rect 221 -737 225 -731
rect 237 -737 241 -731
rect 155 -742 162 -738
rect 166 -742 173 -738
rect 177 -742 184 -738
rect 188 -742 195 -738
rect 151 -748 155 -742
rect 173 -748 177 -742
rect 195 -748 199 -742
rect 161 -771 165 -768
rect 185 -771 189 -768
rect 161 -774 189 -771
rect 129 -781 152 -777
rect 81 -785 85 -781
rect 185 -784 189 -774
rect 230 -784 233 -777
rect 85 -789 91 -785
rect 95 -789 103 -785
rect 107 -789 115 -785
rect 119 -789 125 -785
rect 132 -788 164 -784
rect 185 -788 238 -784
rect 91 -799 98 -795
rect 102 -799 109 -795
rect 113 -799 119 -795
rect 87 -805 91 -799
rect 109 -805 113 -799
rect 75 -838 76 -833
rect 97 -834 101 -825
rect 119 -834 123 -825
rect 81 -838 88 -834
rect 97 -838 123 -834
rect 119 -841 123 -838
rect 132 -841 135 -788
rect 72 -845 100 -841
rect 119 -845 135 -841
rect 138 -795 176 -791
rect 58 -852 112 -848
rect -3 -861 1 -852
rect 23 -861 27 -852
rect -27 -864 -12 -861
rect -3 -865 16 -861
rect -16 -872 0 -869
rect 7 -875 11 -865
rect 23 -866 28 -861
rect 23 -868 27 -866
rect 15 -882 19 -878
rect 19 -886 25 -882
rect 11 -895 57 -892
rect -13 -899 -9 -895
rect -9 -903 -3 -899
rect 1 -903 7 -899
rect 54 -983 57 -895
rect 76 -936 79 -852
rect 119 -855 123 -845
rect 87 -889 91 -885
rect 91 -893 98 -889
rect 102 -893 108 -889
rect 112 -893 119 -889
rect 91 -903 97 -899
rect 101 -903 107 -899
rect 87 -909 91 -903
rect 107 -909 111 -903
rect 75 -938 79 -936
rect 97 -938 101 -929
rect 138 -938 141 -795
rect 75 -941 88 -938
rect 97 -942 141 -938
rect 144 -802 188 -798
rect 78 -949 100 -945
rect 107 -952 111 -942
rect 144 -945 148 -802
rect 195 -805 199 -788
rect 246 -791 249 -777
rect 207 -795 222 -791
rect 226 -795 249 -791
rect 252 -791 255 -731
rect 265 -756 277 -752
rect 261 -762 265 -756
rect 277 -762 281 -756
rect 269 -791 273 -782
rect 285 -791 289 -782
rect 252 -795 262 -791
rect 269 -795 278 -791
rect 285 -795 295 -791
rect 252 -798 255 -795
rect 269 -798 273 -795
rect 285 -798 289 -795
rect 233 -801 255 -798
rect 221 -812 225 -808
rect 261 -812 265 -808
rect 277 -812 281 -808
rect 225 -816 229 -812
rect 233 -816 261 -812
rect 265 -816 269 -812
rect 273 -816 277 -812
rect 281 -816 285 -812
rect 151 -849 155 -845
rect 155 -853 161 -849
rect 165 -853 173 -849
rect 177 -853 185 -849
rect 189 -853 195 -849
rect 114 -948 148 -945
rect 87 -976 91 -972
rect 91 -980 97 -976
rect 101 -980 107 -976
rect 114 -983 117 -948
rect 54 -986 117 -983
rect 79 -998 86 -994
rect 90 -998 97 -994
rect 101 -998 108 -994
rect 112 -998 121 -994
rect 125 -998 131 -994
rect 75 -1004 79 -998
rect 97 -1004 101 -998
rect 121 -1004 125 -998
rect 85 -1027 89 -1024
rect 109 -1027 113 -1024
rect 131 -1027 135 -1024
rect 85 -1030 135 -1027
rect 71 -1037 76 -1033
rect 68 -1042 88 -1040
rect 63 -1044 88 -1042
rect 60 -1051 100 -1047
rect 72 -1058 112 -1054
rect 121 -1062 124 -1051
rect 58 -1065 124 -1062
rect -13 -1112 21 -1108
rect -13 -1118 -9 -1112
rect 3 -1118 7 -1112
rect -4 -1165 -1 -1158
rect -27 -1168 4 -1165
rect -27 -1242 -24 -1168
rect 12 -1172 15 -1158
rect -16 -1176 -12 -1172
rect -8 -1176 15 -1172
rect 18 -1172 21 -1112
rect 31 -1137 43 -1133
rect 27 -1143 31 -1137
rect 43 -1143 47 -1137
rect 35 -1172 39 -1163
rect 51 -1172 55 -1163
rect 58 -1172 61 -1065
rect 131 -1068 135 -1030
rect 135 -1118 141 -1115
rect 75 -1122 79 -1118
rect 79 -1126 85 -1122
rect 89 -1126 97 -1122
rect 101 -1126 109 -1122
rect 113 -1126 121 -1122
rect 125 -1126 131 -1122
rect 87 -1138 94 -1134
rect 98 -1138 105 -1134
rect 109 -1138 116 -1134
rect 120 -1138 127 -1134
rect 83 -1144 87 -1138
rect 105 -1144 109 -1138
rect 127 -1144 131 -1138
rect 93 -1167 97 -1164
rect 117 -1167 121 -1164
rect 93 -1170 121 -1167
rect 18 -1176 28 -1172
rect 35 -1176 44 -1172
rect 51 -1176 61 -1172
rect 18 -1179 21 -1176
rect 35 -1179 39 -1176
rect 51 -1179 55 -1176
rect -1 -1182 21 -1179
rect 58 -1187 61 -1176
rect 78 -1176 84 -1173
rect 117 -1180 121 -1170
rect 138 -1173 141 -1118
rect 158 -1138 165 -1134
rect 169 -1138 176 -1134
rect 180 -1138 187 -1134
rect 191 -1138 200 -1134
rect 204 -1138 210 -1134
rect 154 -1144 158 -1138
rect 176 -1144 180 -1138
rect 200 -1144 204 -1138
rect 164 -1167 168 -1164
rect 188 -1167 192 -1164
rect 210 -1167 214 -1164
rect 164 -1170 214 -1167
rect 138 -1177 155 -1173
rect 69 -1184 96 -1181
rect 117 -1184 167 -1180
rect -13 -1193 -9 -1189
rect 27 -1193 31 -1189
rect 43 -1193 47 -1189
rect 58 -1190 108 -1187
rect -9 -1197 -5 -1193
rect -1 -1197 27 -1193
rect 31 -1197 35 -1193
rect 39 -1197 43 -1193
rect 47 -1197 51 -1193
rect -9 -1207 -3 -1203
rect 1 -1207 7 -1203
rect 11 -1207 15 -1203
rect 19 -1207 25 -1203
rect 29 -1207 33 -1203
rect -13 -1213 -9 -1207
rect 7 -1213 11 -1207
rect 15 -1213 19 -1207
rect -3 -1242 1 -1233
rect -27 -1245 -12 -1242
rect -3 -1246 16 -1242
rect -16 -1253 0 -1250
rect 7 -1256 11 -1246
rect 23 -1249 27 -1233
rect 15 -1263 19 -1259
rect 19 -1267 25 -1263
rect 32 -1272 35 -1256
rect 11 -1276 35 -1272
rect -13 -1280 -9 -1276
rect -9 -1284 -3 -1280
rect 1 -1284 7 -1280
rect 58 -1310 61 -1190
rect 98 -1198 120 -1195
rect 127 -1201 131 -1184
rect 210 -1187 214 -1170
rect 134 -1191 179 -1187
rect 210 -1191 220 -1187
rect 83 -1245 87 -1241
rect 87 -1249 93 -1245
rect 97 -1249 105 -1245
rect 109 -1249 117 -1245
rect 121 -1249 127 -1245
rect 97 -1261 104 -1257
rect 108 -1261 115 -1257
rect 119 -1261 125 -1257
rect 93 -1267 97 -1261
rect 115 -1267 119 -1261
rect 134 -1267 137 -1191
rect 129 -1270 137 -1267
rect 140 -1198 191 -1194
rect 84 -1296 86 -1295
rect 103 -1296 107 -1287
rect 125 -1296 129 -1287
rect 84 -1298 94 -1296
rect 82 -1300 94 -1298
rect 103 -1300 129 -1296
rect 78 -1307 106 -1303
rect 58 -1314 118 -1310
rect 87 -1401 90 -1314
rect 125 -1317 129 -1300
rect 93 -1351 97 -1347
rect 97 -1355 104 -1351
rect 108 -1355 114 -1351
rect 118 -1355 125 -1351
rect 107 -1366 113 -1362
rect 117 -1366 123 -1362
rect 103 -1372 107 -1366
rect 123 -1372 127 -1366
rect 113 -1401 117 -1392
rect 140 -1401 143 -1198
rect 147 -1205 203 -1201
rect 147 -1249 150 -1205
rect 210 -1208 214 -1191
rect 154 -1262 158 -1258
rect 158 -1266 164 -1262
rect 168 -1266 176 -1262
rect 180 -1266 188 -1262
rect 192 -1266 200 -1262
rect 204 -1266 210 -1262
rect 87 -1405 104 -1401
rect 113 -1405 143 -1401
rect 86 -1412 116 -1408
rect 123 -1415 127 -1405
rect 103 -1439 107 -1435
rect 107 -1443 113 -1439
rect 117 -1443 123 -1439
<< m2contact >>
rect 85 -21 90 -16
rect 118 -29 123 -24
rect 53 -43 58 -38
rect -21 -370 -16 -365
rect 93 -378 98 -373
rect -21 -447 -16 -442
rect 30 -470 35 -465
rect 50 -452 55 -447
rect -21 -559 -16 -554
rect 150 -452 155 -447
rect 60 -517 65 -512
rect 50 -581 55 -576
rect -21 -636 -16 -631
rect 23 -630 28 -625
rect -21 -795 -16 -790
rect 74 -724 79 -719
rect 67 -740 72 -735
rect -21 -872 -16 -867
rect 73 -950 78 -945
rect 67 -1059 72 -1054
rect -21 -1176 -16 -1171
rect -21 -1253 -16 -1248
rect 79 -1298 84 -1293
<< metal2 >>
rect 85 -26 89 -21
rect 85 -29 118 -26
rect 85 -43 89 -29
rect 53 -46 89 -43
rect -19 -442 -16 -370
rect 94 -409 97 -378
rect 31 -412 97 -409
rect 31 -465 34 -412
rect 55 -451 150 -448
rect 37 -508 42 -503
rect -19 -631 -16 -559
rect 28 -629 46 -626
rect 43 -744 46 -629
rect 51 -737 54 -581
rect 60 -720 63 -517
rect 67 -574 72 -569
rect 60 -723 74 -720
rect 51 -740 67 -737
rect 43 -747 63 -744
rect -19 -867 -16 -795
rect 60 -945 63 -747
rect 76 -826 79 -724
rect 76 -829 88 -826
rect 85 -851 88 -829
rect 82 -854 88 -851
rect 60 -946 73 -945
rect 41 -949 73 -946
rect 41 -1066 44 -949
rect 82 -987 85 -854
rect 48 -990 85 -987
rect 48 -1055 51 -990
rect 48 -1058 67 -1055
rect 41 -1069 59 -1066
rect -19 -1248 -16 -1176
rect 56 -1294 59 -1069
rect 56 -1298 79 -1294
<< m3contact >>
rect 23 -866 28 -861
<< m123contact >>
rect 132 -349 137 -344
rect 58 -370 63 -365
rect 128 -402 133 -397
rect 129 -444 134 -439
rect 37 -499 42 -494
rect 82 -525 87 -520
rect 67 -614 72 -609
rect 58 -733 63 -728
rect 202 -796 207 -791
rect 76 -838 81 -833
rect 67 -845 72 -840
rect 70 -941 75 -936
rect 70 -1033 75 -1028
rect 63 -1042 68 -1037
rect 55 -1051 60 -1046
rect 120 -1051 125 -1046
rect 31 -1256 36 -1251
rect 73 -1177 78 -1172
rect 64 -1184 69 -1179
rect 93 -1198 98 -1193
rect 146 -1254 151 -1249
rect 73 -1307 78 -1302
rect 81 -1413 86 -1408
<< metal3 >>
rect 128 -349 132 -345
rect 128 -362 131 -349
rect 59 -365 131 -362
rect 38 -503 41 -499
rect 58 -521 61 -370
rect 129 -439 132 -402
rect 58 -525 82 -521
rect 58 -728 61 -525
rect 68 -609 71 -574
rect 28 -865 38 -862
rect 35 -1072 38 -865
rect 59 -920 62 -733
rect 68 -840 71 -614
rect 68 -855 71 -845
rect 56 -923 62 -920
rect 56 -1046 59 -923
rect 78 -928 81 -838
rect 202 -856 205 -796
rect 63 -931 81 -928
rect 151 -859 205 -856
rect 63 -1037 66 -931
rect 70 -1028 73 -941
rect 151 -951 154 -859
rect 140 -954 154 -951
rect 35 -1075 60 -1072
rect 36 -1255 40 -1252
rect 57 -1317 60 -1075
rect 64 -1179 67 -1042
rect 72 -1046 75 -1033
rect 71 -1049 75 -1046
rect 71 -1128 74 -1049
rect 140 -1047 143 -954
rect 125 -1050 143 -1047
rect 71 -1131 76 -1128
rect 73 -1172 76 -1131
rect 73 -1302 76 -1177
rect 85 -1198 93 -1195
rect 85 -1254 146 -1251
rect 57 -1320 84 -1317
rect 81 -1408 84 -1320
<< m345contact >>
rect 37 -508 42 -503
rect 67 -574 72 -569
rect 67 -860 72 -855
rect 80 -1198 85 -1193
rect 40 -1256 45 -1251
rect 80 -1256 85 -1251
<< metal5 >>
rect 42 -507 71 -504
rect 68 -569 71 -507
rect 68 -1195 71 -860
rect 68 -1198 80 -1195
rect 45 -1255 80 -1252
<< labels >>
rlabel metal1 93 -476 93 -476 1 vdd
rlabel metal1 55 -368 55 -368 1 p0
rlabel metal1 123 -368 123 -368 1 c1
rlabel metal1 22 -468 22 -468 1 g0_inv
rlabel metal1 25 -438 25 -438 1 g0
rlabel metal1 118 -329 118 -329 1 vdd
rlabel metal1 68 -375 68 -375 1 c0
rlabel metal1 83 -329 83 -329 1 vdd
rlabel metal1 83 -406 83 -406 1 gnd
rlabel metal2 -18 -373 -18 -373 1 b0
rlabel metal1 -25 -361 -25 -361 1 a0
rlabel metal1 22 -459 22 -459 1 gnd
rlabel metal1 4 -476 4 -476 1 gnd
rlabel metal1 4 -399 4 -399 1 vdd
rlabel metal1 13 -389 13 -389 1 gnd
rlabel metal1 37 -329 37 -329 1 vdd
rlabel metal1 53 -557 53 -557 1 p1
rlabel metal1 22 -648 22 -648 1 gnd
rlabel metal1 4 -665 4 -665 1 gnd
rlabel metal1 4 -588 4 -588 1 vdd
rlabel metal1 13 -578 13 -578 1 gnd
rlabel metal1 37 -518 37 -518 1 vdd
rlabel metal1 -25 -550 -25 -550 1 a1
rlabel metal2 -17 -561 -17 -561 1 b1
rlabel metal1 25 -624 25 -624 1 g1
rlabel metal1 93 -570 93 -570 1 gnd
rlabel metal1 147 -570 147 -570 1 gnd
rlabel metal1 92 -580 92 -580 1 vdd
rlabel metal1 92 -657 92 -657 1 gnd
rlabel metal1 13 -658 13 -658 1 g1_inv
rlabel metal1 -14 -51 -14 -51 1 gnd
rlabel metal1 304 -182 304 -182 7 out_NAND5
rlabel metal1 236 -196 236 -196 1 in5_NAND5
rlabel metal1 236 -189 236 -189 1 in4_NAND5
rlabel metal1 236 -182 236 -182 1 in3_NAND5
rlabel metal1 236 -175 236 -175 1 in2_NAND5
rlabel metal1 236 -168 236 -168 1 in1_NAND5
rlabel metal1 258 -257 258 -257 1 gnd
rlabel metal1 257 -129 257 -129 1 vdd
rlabel space 122 -246 190 -120 1 NAND4
rlabel metal1 184 -175 184 -175 7 out_NAND4
rlabel metal1 128 -189 128 -189 1 in4_NAND4
rlabel metal1 128 -182 128 -182 1 in3_NAND4
rlabel metal1 128 -175 128 -175 1 in2_NAND4
rlabel metal1 128 -168 128 -168 1 in1_NAND4
rlabel metal1 150 -240 150 -240 1 gnd
rlabel metal1 149 -129 149 -129 1 vdd
rlabel space 47 -230 104 -117 1 NAND3
rlabel metal1 98 -175 98 -175 7 out_NAND3
rlabel metal1 76 -223 76 -223 1 gnd
rlabel metal1 76 -129 76 -129 1 vdd
rlabel metal1 54 -182 54 -182 1 in3_NAND3
rlabel metal1 54 -175 54 -175 1 in2_NAND3
rlabel metal1 54 -168 54 -168 1 in1_NAND3
rlabel metal1 15 -168 15 -168 1 out_NAND2
rlabel metal1 4 -206 4 -206 1 gnd
rlabel metal1 -17 -175 -17 -175 1 in2_NAND2
rlabel metal1 -17 -168 -17 -168 1 in1_NAND2
rlabel metal1 4 -129 4 -129 1 vdd
rlabel space -23 -216 28 -119 1 NAND2
rlabel metal1 262 -6 262 -6 1 vdd
rlabel metal1 284 -45 284 -45 1 out_xor
rlabel metal1 208 -45 208 -45 1 in1_xor
rlabel metal1 208 -38 208 -38 1 in2_xor
rlabel space 202 -79 293 29 1 xor
rlabel metal1 238 -66 238 -66 1 gnd
rlabel metal1 -14 9 -14 9 1 vdd
rlabel metal1 -4 -30 -4 -30 1 out_inv
rlabel metal1 -24 -30 -24 -30 1 in_inv
rlabel metal1 170 -21 170 -21 1 out_ff
rlabel metal1 51 -40 51 -40 1 clk
rlabel metal1 51 -49 51 -49 1 in_ff
rlabel space 46 -75 177 26 1 flipflop
rlabel space -33 -60 3 19 1 inverter
rlabel metal1 195 -421 195 -421 5 gnd
rlabel metal1 219 -481 219 -481 5 vdd
rlabel metal1 241 -442 241 -442 1 s1
rlabel metal1 200 -386 200 -386 5 vdd
rlabel metal1 176 -326 176 -326 5 gnd
rlabel metal1 222 -347 222 -347 1 s0
rlabel metal1 218 -1189 218 -1189 1 c4
rlabel metal1 171 -1136 171 -1136 1 vdd
rlabel metal1 172 -1264 172 -1264 1 gnd
rlabel metal1 25 -1244 25 -1244 1 g3
rlabel metal1 13 -1274 13 -1274 1 g3_inv
rlabel metal1 25 -860 25 -860 1 g2
rlabel metal1 120 -1441 120 -1441 1 gnd
rlabel metal1 120 -1364 120 -1364 1 vdd
rlabel metal1 53 -1174 53 -1174 1 p3
rlabel metal1 111 -1353 111 -1353 1 gnd
rlabel metal1 111 -1259 111 -1259 1 vdd
rlabel metal1 101 -1247 101 -1247 1 gnd
rlabel metal1 100 -1136 100 -1136 1 vdd
rlabel metal1 53 -793 53 -793 1 p2
rlabel metal1 93 -1124 93 -1124 1 gnd
rlabel metal1 92 -996 92 -996 1 vdd
rlabel metal1 169 -851 169 -851 1 gnd
rlabel metal1 168 -740 168 -740 1 vdd
rlabel metal1 13 -894 13 -894 1 g2_inv
rlabel metal1 37 -754 37 -754 1 vdd
rlabel metal1 13 -814 13 -814 1 gnd
rlabel metal1 4 -824 4 -824 1 vdd
rlabel metal1 4 -901 4 -901 1 gnd
rlabel metal1 22 -884 22 -884 1 gnd
rlabel metal1 -25 -786 -25 -786 1 a2
rlabel metal2 -17 -797 -17 -797 1 b2
rlabel metal1 98 -676 98 -676 1 vdd
rlabel metal1 99 -787 99 -787 1 gnd
rlabel metal1 105 -797 105 -797 1 vdd
rlabel metal1 105 -891 105 -891 1 gnd
rlabel metal1 104 -978 104 -978 1 gnd
rlabel metal1 104 -901 104 -901 1 vdd
rlabel metal2 -17 -1178 -17 -1178 1 b3
rlabel metal1 -25 -1167 -25 -1167 1 a3
rlabel metal1 37 -1135 37 -1135 1 vdd
rlabel metal1 13 -1195 13 -1195 1 gnd
rlabel metal1 4 -1205 4 -1205 1 vdd
rlabel metal1 4 -1282 4 -1282 1 gnd
rlabel metal1 22 -1265 22 -1265 1 gnd
rlabel metal1 163 -522 163 -522 1 c2
rlabel metal1 177 -648 177 -648 5 gnd
rlabel metal1 201 -708 201 -708 5 vdd
rlabel metal1 224 -669 224 -669 1 s2
rlabel metal1 197 -786 197 -786 1 c3
rlabel metal1 271 -754 271 -754 1 vdd
rlabel metal1 247 -814 247 -814 1 gnd
rlabel metal1 287 -793 287 -793 1 s3
<< end >>
