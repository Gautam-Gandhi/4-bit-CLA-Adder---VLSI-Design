magic
tech scmos
timestamp 1731700802
<< nwell >>
rect -2 -16 22 26
<< ntransistor >>
rect 9 -36 11 -26
<< ptransistor >>
rect 9 -10 11 10
<< ndiffusion >>
rect 8 -36 9 -26
rect 11 -36 12 -26
<< pdiffusion >>
rect 8 -10 9 10
rect 11 -10 12 10
<< ndcontact >>
rect 4 -36 8 -26
rect 12 -36 16 -26
<< pdcontact >>
rect 4 -10 8 10
rect 12 -10 16 10
<< psubstratepcontact >>
rect 0 -46 4 -42
rect 16 -46 20 -42
<< nsubstratencontact >>
rect 1 19 5 23
rect 15 19 19 23
<< polysilicon >>
rect 9 10 11 13
rect 9 -26 11 -10
rect 9 -39 11 -36
<< polycontact >>
rect 5 -23 9 -19
<< metal1 >>
rect -2 23 22 26
rect -2 19 1 23
rect 5 19 15 23
rect 19 19 22 23
rect -2 16 22 19
rect 4 10 8 16
rect 12 -19 16 -10
rect -2 -23 5 -19
rect 12 -23 22 -19
rect 12 -26 16 -23
rect 4 -40 8 -36
rect -2 -42 22 -40
rect -2 -46 0 -42
rect 4 -46 16 -42
rect 20 -46 22 -42
rect -2 -48 22 -46
<< labels >>
rlabel metal1 10 -44 10 -44 1 gnd
rlabel metal1 10 21 10 21 5 vdd
rlabel metal1 0 -21 0 -21 3 in
rlabel metal1 20 -21 20 -21 7 out
<< end >>
