magic
tech scmos
timestamp 1731843905
<< nwell >>
rect -26 -25 -2 14
rect 49 -16 172 23
rect 49 -36 85 -16
rect -32 -109 8 -84
rect -32 -143 48 -109
rect 8 -148 48 -143
<< ntransistor >>
rect -15 -45 -13 -35
rect 96 -50 98 -30
rect 108 -50 110 -30
rect 131 -50 133 -30
rect 143 -50 145 -30
rect 159 -36 161 -26
rect 60 -64 62 -54
rect -21 -168 -19 -158
rect 19 -168 21 -158
rect 35 -168 37 -158
<< ptransistor >>
rect -15 -19 -13 1
rect 60 -30 62 10
rect 72 -30 74 10
rect 96 -10 98 10
rect 131 -10 133 10
rect 159 -10 161 10
rect -21 -137 -19 -97
rect -5 -137 -3 -97
rect 19 -142 21 -122
rect 35 -142 37 -122
<< ndiffusion >>
rect -16 -45 -15 -35
rect -13 -45 -12 -35
rect 95 -50 96 -30
rect 98 -50 108 -30
rect 110 -50 111 -30
rect 130 -50 131 -30
rect 133 -50 143 -30
rect 145 -50 146 -30
rect 158 -36 159 -26
rect 161 -36 162 -26
rect 59 -64 60 -54
rect 62 -64 63 -54
rect -22 -168 -21 -158
rect -19 -168 -18 -158
rect 18 -168 19 -158
rect 21 -168 22 -158
rect 34 -168 35 -158
rect 37 -168 38 -158
<< pdiffusion >>
rect -16 -19 -15 1
rect -13 -19 -12 1
rect 59 -30 60 10
rect 62 -30 72 10
rect 74 -30 75 10
rect 95 -10 96 10
rect 98 -10 99 10
rect 130 -10 131 10
rect 133 -10 134 10
rect 158 -10 159 10
rect 161 -10 162 10
rect -22 -137 -21 -97
rect -19 -137 -18 -97
rect -6 -137 -5 -97
rect -3 -137 -2 -97
rect 18 -142 19 -122
rect 21 -142 22 -122
rect 34 -142 35 -122
rect 37 -142 38 -122
<< ndcontact >>
rect -20 -45 -16 -35
rect -12 -45 -8 -35
rect 91 -50 95 -30
rect 111 -50 115 -30
rect 126 -50 130 -30
rect 146 -50 150 -30
rect 154 -36 158 -26
rect 162 -36 166 -26
rect 55 -64 59 -54
rect 63 -64 67 -54
rect -26 -168 -22 -158
rect -18 -168 -14 -158
rect 14 -168 18 -158
rect 22 -168 26 -158
rect 30 -168 34 -158
rect 38 -168 42 -158
<< pdcontact >>
rect -20 -19 -16 1
rect -12 -19 -8 1
rect 55 -30 59 10
rect 75 -30 79 10
rect 91 -10 95 10
rect 99 -10 103 10
rect 126 -10 130 10
rect 134 -10 138 10
rect 154 -10 158 10
rect 162 -10 166 10
rect -26 -137 -22 -97
rect -18 -137 -14 -97
rect -10 -137 -6 -97
rect -2 -137 2 -97
rect 14 -142 18 -122
rect 22 -142 26 -122
rect 30 -142 34 -122
rect 38 -142 42 -122
<< psubstratepcontact >>
rect -20 -53 -16 -49
rect -10 -53 -6 -49
rect 154 -44 158 -40
rect 164 -44 168 -40
rect 72 -58 76 -54
rect 87 -58 91 -54
rect 103 -58 107 -54
rect 122 -58 126 -54
rect 138 -58 142 -54
rect 154 -58 158 -54
rect 51 -72 55 -68
rect 62 -72 66 -68
rect 72 -72 76 -68
rect -26 -176 -22 -172
rect -18 -176 -14 -172
rect 14 -176 18 -172
rect 22 -176 26 -172
rect 30 -176 34 -172
rect 38 -176 42 -172
<< nsubstratencontact >>
rect 53 16 57 20
rect 65 16 69 20
rect 76 16 80 20
rect 87 16 91 20
rect 101 16 105 20
rect 112 16 116 20
rect 122 16 126 20
rect 136 16 140 20
rect 152 16 156 20
rect 164 16 168 20
rect -22 7 -18 11
rect -10 7 -6 11
rect 14 -116 18 -112
rect 30 -116 34 -112
<< polysilicon >>
rect 60 10 62 13
rect 72 10 74 13
rect 96 10 98 13
rect 131 10 133 13
rect 159 10 161 13
rect -15 1 -13 4
rect -15 -35 -13 -19
rect 96 -30 98 -10
rect 108 -30 110 -23
rect 131 -30 133 -10
rect 143 -30 145 -23
rect 159 -26 161 -10
rect -15 -48 -13 -45
rect 60 -54 62 -30
rect 72 -44 74 -30
rect 159 -39 161 -36
rect 96 -53 98 -50
rect 108 -53 110 -50
rect 131 -53 133 -50
rect 143 -53 145 -50
rect 60 -67 62 -64
rect -21 -97 -19 -94
rect -5 -97 -3 -94
rect 19 -122 21 -119
rect 35 -122 37 -119
rect -21 -158 -19 -137
rect -5 -148 -3 -137
rect 19 -158 21 -142
rect 35 -158 37 -142
rect -21 -171 -19 -168
rect 19 -171 21 -168
rect 35 -171 37 -168
<< polycontact >>
rect -19 -32 -15 -28
rect 92 -20 96 -16
rect 127 -21 131 -17
rect 104 -27 108 -23
rect 155 -23 159 -19
rect 139 -27 143 -23
rect 56 -51 60 -47
rect 68 -42 72 -38
rect -25 -155 -21 -151
rect -9 -148 -5 -144
rect 15 -155 19 -151
rect 31 -155 35 -151
<< metal1 >>
rect 49 16 53 20
rect 57 16 65 20
rect 69 16 76 20
rect 80 16 87 20
rect 91 16 101 20
rect 105 16 112 20
rect 116 16 122 20
rect 126 16 136 20
rect 140 16 152 20
rect 156 16 164 20
rect 168 16 172 20
rect -26 7 -22 11
rect -18 7 -10 11
rect -6 7 -2 11
rect 55 10 59 16
rect 91 10 95 16
rect 126 10 130 16
rect 154 10 158 16
rect -20 1 -16 7
rect -12 -28 -8 -19
rect -26 -32 -19 -28
rect -12 -32 -2 -28
rect 90 -20 92 -16
rect 99 -17 103 -10
rect 134 -17 138 -10
rect 99 -20 127 -17
rect 111 -21 127 -20
rect 134 -19 150 -17
rect 162 -19 166 -10
rect 134 -20 155 -19
rect 79 -27 104 -24
rect 111 -30 115 -21
rect 146 -23 155 -20
rect 162 -23 172 -19
rect 123 -27 139 -24
rect 146 -30 150 -23
rect 162 -26 166 -23
rect -12 -35 -8 -32
rect 49 -42 53 -38
rect 58 -42 68 -38
rect -20 -49 -16 -45
rect 75 -47 79 -30
rect -26 -53 -20 -49
rect -16 -53 -10 -49
rect -6 -53 -2 -49
rect 49 -51 56 -47
rect 63 -51 79 -47
rect 154 -40 158 -36
rect 158 -44 164 -40
rect 168 -44 172 -40
rect 63 -54 67 -51
rect 91 -54 95 -50
rect 126 -54 130 -50
rect 154 -54 158 -44
rect 76 -58 87 -54
rect 91 -58 103 -54
rect 107 -58 122 -54
rect 126 -58 138 -54
rect 142 -58 154 -54
rect 55 -68 59 -64
rect 72 -68 76 -58
rect 49 -72 51 -68
rect 55 -72 62 -68
rect 66 -72 72 -68
rect -32 -91 8 -87
rect -26 -97 -22 -91
rect -10 -97 -6 -91
rect -17 -144 -14 -137
rect -32 -148 -9 -144
rect -1 -151 2 -137
rect -32 -155 -25 -151
rect -21 -155 2 -151
rect 5 -151 8 -91
rect 18 -116 30 -112
rect 14 -122 18 -116
rect 30 -122 34 -116
rect 22 -151 26 -142
rect 38 -151 42 -142
rect 5 -155 15 -151
rect 22 -155 31 -151
rect 38 -155 48 -151
rect 5 -158 8 -155
rect 22 -158 26 -155
rect 38 -158 42 -155
rect -14 -161 8 -158
rect -26 -172 -22 -168
rect 14 -172 18 -168
rect 30 -172 34 -168
rect -32 -176 -26 -172
rect -22 -176 -18 -172
rect -14 -176 14 -172
rect 18 -176 22 -172
rect 26 -176 30 -172
rect 34 -176 38 -172
<< m2contact >>
rect 85 -21 90 -16
rect 118 -29 123 -24
rect 53 -43 58 -38
<< metal2 >>
rect 85 -26 89 -21
rect 85 -29 118 -26
rect 85 -43 89 -29
rect 53 -46 89 -43
<< labels >>
rlabel space -33 -60 3 19 1 inverter
rlabel space 46 -75 177 26 1 flipflop
rlabel metal1 -30 -153 -30 -153 3 in1
rlabel metal1 -30 -146 -30 -146 3 in2
rlabel metal1 0 -174 0 -174 1 gnd
rlabel metal1 51 -49 51 -49 1 in_ff
rlabel metal1 51 -40 51 -40 1 clk
rlabel metal1 170 -21 170 -21 1 out_ff
rlabel metal1 24 -114 24 -114 1 vdd
rlabel metal1 -24 -30 -24 -30 1 in_inv
rlabel metal1 -4 -30 -4 -30 1 out_inv
rlabel metal1 -14 9 -14 9 1 vdd
rlabel metal1 -13 -51 -13 -51 1 gnd
rlabel metal1 46 -153 46 -153 1 out_xor
<< end >>
